module RGB2GrayFilter(
  input         clock,
  input         reset,
  output        io_enq_ready,
  input         io_enq_valid,
  input  [23:0] io_enq_bits,
  input         io_enq_user,
  input         io_enq_last,
  input         io_deq_ready,
  output        io_deq_valid,
  output [23:0] io_deq_bits,
  output        io_deq_user,
  output        io_deq_last,
  output [8:0]  xcounter_0,
  output [8:0]  ycounter_0
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
`endif // RANDOMIZE_REG_INIT
  reg [1:0] stateReg; // @[ChiselImProc.scala 62:28]
  reg [23:0] dataReg; // @[ChiselImProc.scala 64:23]
  reg [23:0] shadowReg; // @[ChiselImProc.scala 66:25]
  reg  userReg; // @[ChiselImProc.scala 67:23]
  reg  shadowUserReg; // @[ChiselImProc.scala 68:29]
  reg  lastReg; // @[ChiselImProc.scala 69:23]
  reg  shadowLastReg; // @[ChiselImProc.scala 70:29]
  wire  _T = 2'h0 == stateReg; // @[Conditional.scala 37:30]
  wire  _T_1 = 2'h1 == stateReg; // @[Conditional.scala 37:30]
  wire  _T_2 = ~io_enq_valid; // @[ChiselImProc.scala 84:39]
  wire  _T_3 = io_deq_ready & _T_2; // @[ChiselImProc.scala 84:36]
  wire  _T_4 = io_deq_ready & io_enq_valid; // @[ChiselImProc.scala 87:42]
  wire  _T_5 = ~io_deq_ready; // @[ChiselImProc.scala 92:29]
  wire  _T_6 = _T_5 & io_enq_valid; // @[ChiselImProc.scala 92:43]
  wire  _T_7 = 2'h2 == stateReg; // @[Conditional.scala 37:30]
  wire  _T_8 = 2'h3 == stateReg; // @[Conditional.scala 37:30]
  wire  _T_9 = stateReg == 2'h0; // @[ChiselImProc.scala 116:35]
  wire  _T_10 = stateReg == 2'h1; // @[ChiselImProc.scala 116:57]
  wire  _T_11 = _T_9 | _T_10; // @[ChiselImProc.scala 116:45]
  wire  _T_12 = stateReg == 2'h3; // @[ChiselImProc.scala 116:77]
  wire  _T_15 = stateReg == 2'h2; // @[ChiselImProc.scala 117:55]
  wire  _T_16 = _T_10 | _T_15; // @[ChiselImProc.scala 117:43]
  reg [8:0] xcounter; // @[ChiselImProc.scala 170:23]
  reg [8:0] ycounter; // @[ChiselImProc.scala 171:23]
  wire  _T_20 = lastReg & _T_16; // @[ChiselImProc.scala 176:25]
  wire  _T_21 = _T_20 & io_deq_ready; // @[ChiselImProc.scala 176:67]
  wire [8:0] _T_23 = ycounter + 9'h1; // @[ChiselImProc.scala 178:30]
  wire  _T_27 = _T_16 & io_deq_ready; // @[ChiselImProc.scala 179:56]
  wire [8:0] _T_29 = xcounter + 9'h1; // @[ChiselImProc.scala 180:30]
  wire [23:0] _T_30 = dataReg & 24'hff; // @[ChiselImProc.scala 186:36]
  wire [37:0] _T_31 = 24'h24dd * _T_30; // @[ChiselImProc.scala 186:25]
  wire [23:0] _T_32 = dataReg & 24'hff00; // @[ChiselImProc.scala 187:33]
  wire [23:0] _T_33 = {{8'd0}, _T_32[23:8]}; // @[ChiselImProc.scala 187:47]
  wire [39:0] _T_34 = 24'h9645 * _T_33; // @[ChiselImProc.scala 187:21]
  wire [39:0] _GEN_50 = {{2'd0}, _T_31}; // @[ChiselImProc.scala 186:50]
  wire [39:0] _T_36 = _GEN_50 + _T_34; // @[ChiselImProc.scala 186:50]
  wire [23:0] _T_37 = dataReg & 24'hff0000; // @[ChiselImProc.scala 188:33]
  wire [23:0] _T_38 = {{16'd0}, _T_37[23:16]}; // @[ChiselImProc.scala 188:47]
  wire [38:0] _T_39 = 24'h4c8b * _T_38; // @[ChiselImProc.scala 188:21]
  wire [39:0] _GEN_52 = {{1'd0}, _T_39}; // @[ChiselImProc.scala 187:55]
  wire [39:0] _T_41 = _T_36 + _GEN_52; // @[ChiselImProc.scala 187:55]
  wire [31:0] pixGray = _T_41[31:0]; // @[ChiselImProc.scala 166:24 ChiselImProc.scala 186:13]
  wire [31:0] _T_42 = {{16'd0}, pixGray[31:16]}; // @[ChiselImProc.scala 190:24]
  wire [15:0] rolled = _T_42[15:0]; // @[ChiselImProc.scala 167:23 ChiselImProc.scala 190:12]
  wire  _T_43 = rolled > 16'hff; // @[ChiselImProc.scala 191:32]
  wire [15:0] _T_44 = _T_43 ? 16'hff : rolled; // @[ChiselImProc.scala 191:24]
  assign io_enq_ready = _T_11 | _T_12; // @[ChiselImProc.scala 116:22]
  assign io_deq_valid = _T_10 | _T_15; // @[ChiselImProc.scala 117:22]
  assign io_deq_bits = {{8'd0}, _T_44}; // @[ChiselImProc.scala 191:17]
  assign io_deq_user = userReg; // @[ChiselImProc.scala 144:17 ChiselImProc.scala 114:21]
  assign io_deq_last = lastReg; // @[ChiselImProc.scala 143:17 ChiselImProc.scala 113:21]
  assign xcounter_0 = xcounter;
  assign ycounter_0 = ycounter;
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  stateReg = _RAND_0[1:0];
  _RAND_1 = {1{`RANDOM}};
  dataReg = _RAND_1[23:0];
  _RAND_2 = {1{`RANDOM}};
  shadowReg = _RAND_2[23:0];
  _RAND_3 = {1{`RANDOM}};
  userReg = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  shadowUserReg = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  lastReg = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  shadowLastReg = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  xcounter = _RAND_7[8:0];
  _RAND_8 = {1{`RANDOM}};
  ycounter = _RAND_8[8:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      stateReg <= 2'h0;
    end else if (_T) begin
      if (io_enq_valid) begin
        stateReg <= 2'h1;
      end
    end else if (_T_1) begin
      if (_T_3) begin
        stateReg <= 2'h0;
      end else if (_T_4) begin
        stateReg <= 2'h1;
      end else if (_T_6) begin
        stateReg <= 2'h2;
      end
    end else if (_T_7) begin
      if (io_deq_ready) begin
        stateReg <= 2'h1;
      end
    end else if (_T_8) begin
      stateReg <= 2'h0;
    end
    if (_T) begin
      if (io_enq_valid) begin
        dataReg <= io_enq_bits;
      end
    end else if (_T_1) begin
      if (!(_T_3)) begin
        if (_T_4) begin
          dataReg <= io_enq_bits;
        end
      end
    end else if (_T_7) begin
      if (io_deq_ready) begin
        dataReg <= shadowReg;
      end
    end
    if (!(_T)) begin
      if (_T_1) begin
        if (!(_T_3)) begin
          if (!(_T_4)) begin
            if (_T_6) begin
              shadowReg <= io_enq_bits;
            end
          end
        end
      end
    end
    if (_T) begin
      userReg <= io_enq_user;
    end else if (_T_1) begin
      if (_T_3) begin
        userReg <= io_enq_user;
      end else if (_T_4) begin
        userReg <= io_enq_user;
      end
    end else if (_T_7) begin
      if (io_deq_ready) begin
        userReg <= shadowUserReg;
      end
    end
    if (!(_T)) begin
      if (_T_1) begin
        if (!(_T_3)) begin
          if (!(_T_4)) begin
            if (_T_6) begin
              shadowUserReg <= io_enq_user;
            end
          end
        end
      end
    end
    if (_T) begin
      if (io_enq_valid) begin
        lastReg <= io_enq_last;
      end
    end else if (_T_1) begin
      if (!(_T_3)) begin
        if (_T_4) begin
          lastReg <= io_enq_last;
        end
      end
    end else if (_T_7) begin
      if (io_deq_ready) begin
        lastReg <= shadowLastReg;
      end
    end
    if (!(_T)) begin
      if (_T_1) begin
        if (!(_T_3)) begin
          if (!(_T_4)) begin
            if (_T_6) begin
              shadowLastReg <= io_enq_last;
            end
          end
        end
      end
    end
    if (userReg) begin
      xcounter <= 9'h0;
    end else if (_T_21) begin
      xcounter <= 9'h0;
    end else if (_T_27) begin
      xcounter <= _T_29;
    end
    if (userReg) begin
      ycounter <= 9'h0;
    end else if (_T_21) begin
      ycounter <= _T_23;
    end
  end
endmodule
module MulAdd(
  input  [7:0]  io__b_0,
  input  [7:0]  io__b_1,
  input  [7:0]  io__b_2,
  input  [7:0]  io__b_3,
  input  [7:0]  io__b_4,
  input  [7:0]  io__b_5,
  input  [7:0]  io__b_6,
  input  [7:0]  io__b_7,
  input  [7:0]  io__b_8,
  output [15:0] io__output,
  output [15:0] io_output
);
  wire [15:0] _T = 8'h1 * io__b_0; // @[ChiselImProc.scala 32:32]
  wire [16:0] _T_1 = {{1'd0}, _T}; // @[ChiselImProc.scala 32:19]
  wire [15:0] _T_3 = 8'h2 * io__b_1; // @[ChiselImProc.scala 32:32]
  wire [15:0] _T_5 = _T_1[15:0] + _T_3; // @[ChiselImProc.scala 32:19]
  wire [15:0] _T_6 = 8'h1 * io__b_2; // @[ChiselImProc.scala 32:32]
  wire [15:0] _T_8 = _T_5 + _T_6; // @[ChiselImProc.scala 32:19]
  wire [16:0] _T_9 = {{1'd0}, _T_8}; // @[ChiselImProc.scala 34:13]
  wire [15:0] _T_11 = 8'h2 * io__b_3; // @[ChiselImProc.scala 32:32]
  wire [16:0] _T_12 = {{1'd0}, _T_11}; // @[ChiselImProc.scala 32:19]
  wire [15:0] _T_14 = 8'h4 * io__b_4; // @[ChiselImProc.scala 32:32]
  wire [15:0] _T_16 = _T_12[15:0] + _T_14; // @[ChiselImProc.scala 32:19]
  wire [15:0] _T_17 = 8'h2 * io__b_5; // @[ChiselImProc.scala 32:32]
  wire [15:0] _T_19 = _T_16 + _T_17; // @[ChiselImProc.scala 32:19]
  wire [15:0] _T_21 = _T_9[15:0] + _T_19; // @[ChiselImProc.scala 34:13]
  wire [15:0] _T_22 = 8'h1 * io__b_6; // @[ChiselImProc.scala 32:32]
  wire [16:0] _T_23 = {{1'd0}, _T_22}; // @[ChiselImProc.scala 32:19]
  wire [15:0] _T_25 = 8'h2 * io__b_7; // @[ChiselImProc.scala 32:32]
  wire [15:0] _T_27 = _T_23[15:0] + _T_25; // @[ChiselImProc.scala 32:19]
  wire [15:0] _T_28 = 8'h1 * io__b_8; // @[ChiselImProc.scala 32:32]
  wire [15:0] _T_30 = _T_27 + _T_28; // @[ChiselImProc.scala 32:19]
  assign io__output = _T_21 + _T_30; // @[ChiselImProc.scala 36:15]
  assign io_output = io__output;
endmodule
module GaussianBlurFilter(
  input         clock,
  input         reset,
  output        io__enq_ready,
  input         io__enq_valid,
  input  [7:0]  io__enq_bits,
  input         io__enq_user,
  input         io__enq_last,
  input         io__deq_ready,
  output        io__deq_valid,
  output [7:0]  io__deq_bits,
  output        io__deq_user,
  output        io__deq_last,
  output        io_deq_ready,
  output        io_deq_valid,
  output [71:0] _T_805_0,
  output [15:0] io_output
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
  reg [31:0] _RAND_64;
  reg [31:0] _RAND_65;
  reg [31:0] _RAND_66;
  reg [31:0] _RAND_67;
  reg [31:0] _RAND_68;
  reg [31:0] _RAND_69;
  reg [31:0] _RAND_70;
  reg [31:0] _RAND_71;
  reg [31:0] _RAND_72;
  reg [31:0] _RAND_73;
  reg [31:0] _RAND_74;
  reg [31:0] _RAND_75;
  reg [31:0] _RAND_76;
  reg [31:0] _RAND_77;
  reg [31:0] _RAND_78;
  reg [31:0] _RAND_79;
  reg [31:0] _RAND_80;
  reg [31:0] _RAND_81;
  reg [31:0] _RAND_82;
  reg [31:0] _RAND_83;
  reg [31:0] _RAND_84;
  reg [31:0] _RAND_85;
  reg [31:0] _RAND_86;
  reg [31:0] _RAND_87;
  reg [31:0] _RAND_88;
  reg [31:0] _RAND_89;
  reg [31:0] _RAND_90;
  reg [31:0] _RAND_91;
  reg [31:0] _RAND_92;
  reg [31:0] _RAND_93;
  reg [31:0] _RAND_94;
  reg [31:0] _RAND_95;
  reg [31:0] _RAND_96;
  reg [31:0] _RAND_97;
  reg [31:0] _RAND_98;
  reg [31:0] _RAND_99;
  reg [31:0] _RAND_100;
  reg [31:0] _RAND_101;
  reg [31:0] _RAND_102;
  reg [31:0] _RAND_103;
  reg [31:0] _RAND_104;
  reg [31:0] _RAND_105;
  reg [31:0] _RAND_106;
  reg [31:0] _RAND_107;
  reg [31:0] _RAND_108;
  reg [31:0] _RAND_109;
  reg [31:0] _RAND_110;
  reg [31:0] _RAND_111;
  reg [31:0] _RAND_112;
  reg [31:0] _RAND_113;
  reg [31:0] _RAND_114;
  reg [31:0] _RAND_115;
  reg [31:0] _RAND_116;
  reg [31:0] _RAND_117;
  reg [31:0] _RAND_118;
  reg [31:0] _RAND_119;
  reg [31:0] _RAND_120;
  reg [31:0] _RAND_121;
  reg [31:0] _RAND_122;
  reg [31:0] _RAND_123;
  reg [31:0] _RAND_124;
  reg [31:0] _RAND_125;
  reg [31:0] _RAND_126;
  reg [31:0] _RAND_127;
  reg [31:0] _RAND_128;
  reg [31:0] _RAND_129;
  reg [31:0] _RAND_130;
  reg [31:0] _RAND_131;
  reg [31:0] _RAND_132;
  reg [31:0] _RAND_133;
  reg [31:0] _RAND_134;
  reg [31:0] _RAND_135;
  reg [31:0] _RAND_136;
  reg [31:0] _RAND_137;
  reg [31:0] _RAND_138;
  reg [31:0] _RAND_139;
  reg [31:0] _RAND_140;
  reg [31:0] _RAND_141;
  reg [31:0] _RAND_142;
  reg [31:0] _RAND_143;
  reg [31:0] _RAND_144;
  reg [31:0] _RAND_145;
  reg [31:0] _RAND_146;
  reg [31:0] _RAND_147;
  reg [31:0] _RAND_148;
  reg [31:0] _RAND_149;
  reg [31:0] _RAND_150;
  reg [31:0] _RAND_151;
  reg [31:0] _RAND_152;
  reg [31:0] _RAND_153;
  reg [31:0] _RAND_154;
  reg [31:0] _RAND_155;
  reg [31:0] _RAND_156;
  reg [31:0] _RAND_157;
  reg [31:0] _RAND_158;
  reg [31:0] _RAND_159;
  reg [31:0] _RAND_160;
  reg [31:0] _RAND_161;
  reg [31:0] _RAND_162;
  reg [31:0] _RAND_163;
  reg [31:0] _RAND_164;
  reg [31:0] _RAND_165;
  reg [31:0] _RAND_166;
  reg [31:0] _RAND_167;
  reg [31:0] _RAND_168;
  reg [31:0] _RAND_169;
  reg [31:0] _RAND_170;
  reg [31:0] _RAND_171;
  reg [31:0] _RAND_172;
  reg [31:0] _RAND_173;
  reg [31:0] _RAND_174;
  reg [31:0] _RAND_175;
  reg [31:0] _RAND_176;
  reg [31:0] _RAND_177;
  reg [31:0] _RAND_178;
  reg [31:0] _RAND_179;
  reg [31:0] _RAND_180;
  reg [31:0] _RAND_181;
  reg [31:0] _RAND_182;
  reg [31:0] _RAND_183;
  reg [31:0] _RAND_184;
  reg [31:0] _RAND_185;
  reg [31:0] _RAND_186;
  reg [31:0] _RAND_187;
  reg [31:0] _RAND_188;
  reg [31:0] _RAND_189;
  reg [31:0] _RAND_190;
  reg [31:0] _RAND_191;
  reg [31:0] _RAND_192;
  reg [31:0] _RAND_193;
  reg [31:0] _RAND_194;
  reg [31:0] _RAND_195;
  reg [31:0] _RAND_196;
  reg [31:0] _RAND_197;
  reg [31:0] _RAND_198;
  reg [31:0] _RAND_199;
  reg [31:0] _RAND_200;
  reg [31:0] _RAND_201;
  reg [31:0] _RAND_202;
  reg [31:0] _RAND_203;
  reg [31:0] _RAND_204;
  reg [31:0] _RAND_205;
  reg [31:0] _RAND_206;
  reg [31:0] _RAND_207;
  reg [31:0] _RAND_208;
  reg [31:0] _RAND_209;
  reg [31:0] _RAND_210;
  reg [31:0] _RAND_211;
  reg [31:0] _RAND_212;
  reg [31:0] _RAND_213;
  reg [31:0] _RAND_214;
  reg [31:0] _RAND_215;
  reg [31:0] _RAND_216;
  reg [31:0] _RAND_217;
  reg [31:0] _RAND_218;
  reg [31:0] _RAND_219;
  reg [31:0] _RAND_220;
  reg [31:0] _RAND_221;
  reg [31:0] _RAND_222;
  reg [31:0] _RAND_223;
  reg [31:0] _RAND_224;
  reg [31:0] _RAND_225;
  reg [31:0] _RAND_226;
  reg [31:0] _RAND_227;
  reg [31:0] _RAND_228;
  reg [31:0] _RAND_229;
  reg [31:0] _RAND_230;
  reg [31:0] _RAND_231;
  reg [31:0] _RAND_232;
  reg [31:0] _RAND_233;
  reg [31:0] _RAND_234;
  reg [31:0] _RAND_235;
  reg [31:0] _RAND_236;
  reg [31:0] _RAND_237;
  reg [31:0] _RAND_238;
  reg [31:0] _RAND_239;
  reg [31:0] _RAND_240;
  reg [31:0] _RAND_241;
  reg [31:0] _RAND_242;
  reg [31:0] _RAND_243;
  reg [31:0] _RAND_244;
  reg [31:0] _RAND_245;
  reg [31:0] _RAND_246;
  reg [31:0] _RAND_247;
  reg [31:0] _RAND_248;
  reg [31:0] _RAND_249;
  reg [31:0] _RAND_250;
  reg [31:0] _RAND_251;
  reg [31:0] _RAND_252;
  reg [31:0] _RAND_253;
  reg [31:0] _RAND_254;
  reg [31:0] _RAND_255;
  reg [31:0] _RAND_256;
  reg [31:0] _RAND_257;
  reg [31:0] _RAND_258;
  reg [31:0] _RAND_259;
  reg [31:0] _RAND_260;
  reg [31:0] _RAND_261;
  reg [31:0] _RAND_262;
  reg [31:0] _RAND_263;
  reg [31:0] _RAND_264;
  reg [31:0] _RAND_265;
  reg [31:0] _RAND_266;
  reg [31:0] _RAND_267;
  reg [31:0] _RAND_268;
  reg [31:0] _RAND_269;
  reg [31:0] _RAND_270;
  reg [31:0] _RAND_271;
  reg [31:0] _RAND_272;
  reg [31:0] _RAND_273;
  reg [31:0] _RAND_274;
  reg [31:0] _RAND_275;
  reg [31:0] _RAND_276;
  reg [31:0] _RAND_277;
  reg [31:0] _RAND_278;
  reg [31:0] _RAND_279;
  reg [31:0] _RAND_280;
  reg [31:0] _RAND_281;
  reg [31:0] _RAND_282;
  reg [31:0] _RAND_283;
  reg [31:0] _RAND_284;
  reg [31:0] _RAND_285;
  reg [31:0] _RAND_286;
  reg [31:0] _RAND_287;
  reg [31:0] _RAND_288;
  reg [31:0] _RAND_289;
  reg [31:0] _RAND_290;
  reg [31:0] _RAND_291;
  reg [31:0] _RAND_292;
  reg [31:0] _RAND_293;
  reg [31:0] _RAND_294;
  reg [31:0] _RAND_295;
  reg [31:0] _RAND_296;
  reg [31:0] _RAND_297;
  reg [31:0] _RAND_298;
  reg [31:0] _RAND_299;
  reg [31:0] _RAND_300;
  reg [31:0] _RAND_301;
  reg [31:0] _RAND_302;
  reg [31:0] _RAND_303;
  reg [31:0] _RAND_304;
  reg [31:0] _RAND_305;
  reg [31:0] _RAND_306;
  reg [31:0] _RAND_307;
  reg [31:0] _RAND_308;
  reg [31:0] _RAND_309;
  reg [31:0] _RAND_310;
  reg [31:0] _RAND_311;
  reg [31:0] _RAND_312;
  reg [31:0] _RAND_313;
  reg [31:0] _RAND_314;
  reg [31:0] _RAND_315;
  reg [31:0] _RAND_316;
  reg [31:0] _RAND_317;
  reg [31:0] _RAND_318;
  reg [31:0] _RAND_319;
  reg [31:0] _RAND_320;
  reg [31:0] _RAND_321;
  reg [31:0] _RAND_322;
  reg [31:0] _RAND_323;
  reg [31:0] _RAND_324;
  reg [31:0] _RAND_325;
  reg [31:0] _RAND_326;
  reg [31:0] _RAND_327;
  reg [31:0] _RAND_328;
  reg [31:0] _RAND_329;
  reg [31:0] _RAND_330;
  reg [31:0] _RAND_331;
  reg [31:0] _RAND_332;
  reg [31:0] _RAND_333;
  reg [31:0] _RAND_334;
  reg [31:0] _RAND_335;
  reg [31:0] _RAND_336;
  reg [31:0] _RAND_337;
  reg [31:0] _RAND_338;
  reg [31:0] _RAND_339;
  reg [31:0] _RAND_340;
  reg [31:0] _RAND_341;
  reg [31:0] _RAND_342;
  reg [31:0] _RAND_343;
  reg [31:0] _RAND_344;
  reg [31:0] _RAND_345;
  reg [31:0] _RAND_346;
  reg [31:0] _RAND_347;
  reg [31:0] _RAND_348;
  reg [31:0] _RAND_349;
  reg [31:0] _RAND_350;
  reg [31:0] _RAND_351;
  reg [31:0] _RAND_352;
  reg [31:0] _RAND_353;
  reg [31:0] _RAND_354;
  reg [31:0] _RAND_355;
  reg [31:0] _RAND_356;
  reg [31:0] _RAND_357;
  reg [31:0] _RAND_358;
  reg [31:0] _RAND_359;
  reg [31:0] _RAND_360;
  reg [31:0] _RAND_361;
  reg [31:0] _RAND_362;
  reg [31:0] _RAND_363;
  reg [31:0] _RAND_364;
  reg [31:0] _RAND_365;
  reg [31:0] _RAND_366;
  reg [31:0] _RAND_367;
  reg [31:0] _RAND_368;
  reg [31:0] _RAND_369;
  reg [31:0] _RAND_370;
  reg [31:0] _RAND_371;
  reg [31:0] _RAND_372;
  reg [31:0] _RAND_373;
  reg [31:0] _RAND_374;
  reg [31:0] _RAND_375;
  reg [31:0] _RAND_376;
  reg [31:0] _RAND_377;
  reg [31:0] _RAND_378;
  reg [31:0] _RAND_379;
  reg [31:0] _RAND_380;
  reg [31:0] _RAND_381;
  reg [31:0] _RAND_382;
  reg [31:0] _RAND_383;
  reg [31:0] _RAND_384;
  reg [31:0] _RAND_385;
  reg [31:0] _RAND_386;
  reg [31:0] _RAND_387;
  reg [31:0] _RAND_388;
  reg [31:0] _RAND_389;
  reg [31:0] _RAND_390;
  reg [31:0] _RAND_391;
  reg [31:0] _RAND_392;
  reg [31:0] _RAND_393;
  reg [31:0] _RAND_394;
  reg [31:0] _RAND_395;
  reg [31:0] _RAND_396;
  reg [31:0] _RAND_397;
  reg [31:0] _RAND_398;
  reg [31:0] _RAND_399;
  reg [31:0] _RAND_400;
  reg [31:0] _RAND_401;
  reg [31:0] _RAND_402;
  reg [31:0] _RAND_403;
  reg [31:0] _RAND_404;
  reg [31:0] _RAND_405;
  reg [31:0] _RAND_406;
  reg [31:0] _RAND_407;
  reg [31:0] _RAND_408;
  reg [31:0] _RAND_409;
  reg [31:0] _RAND_410;
  reg [31:0] _RAND_411;
  reg [31:0] _RAND_412;
  reg [31:0] _RAND_413;
  reg [31:0] _RAND_414;
  reg [31:0] _RAND_415;
  reg [31:0] _RAND_416;
  reg [31:0] _RAND_417;
  reg [31:0] _RAND_418;
  reg [31:0] _RAND_419;
  reg [31:0] _RAND_420;
  reg [31:0] _RAND_421;
  reg [31:0] _RAND_422;
  reg [31:0] _RAND_423;
  reg [31:0] _RAND_424;
  reg [31:0] _RAND_425;
  reg [31:0] _RAND_426;
  reg [31:0] _RAND_427;
  reg [31:0] _RAND_428;
  reg [31:0] _RAND_429;
  reg [31:0] _RAND_430;
  reg [31:0] _RAND_431;
  reg [31:0] _RAND_432;
  reg [31:0] _RAND_433;
  reg [31:0] _RAND_434;
  reg [31:0] _RAND_435;
  reg [31:0] _RAND_436;
  reg [31:0] _RAND_437;
  reg [31:0] _RAND_438;
  reg [31:0] _RAND_439;
  reg [31:0] _RAND_440;
  reg [31:0] _RAND_441;
  reg [31:0] _RAND_442;
  reg [31:0] _RAND_443;
  reg [31:0] _RAND_444;
  reg [31:0] _RAND_445;
  reg [31:0] _RAND_446;
  reg [31:0] _RAND_447;
  reg [31:0] _RAND_448;
  reg [31:0] _RAND_449;
  reg [31:0] _RAND_450;
  reg [31:0] _RAND_451;
  reg [31:0] _RAND_452;
  reg [31:0] _RAND_453;
  reg [31:0] _RAND_454;
  reg [31:0] _RAND_455;
  reg [31:0] _RAND_456;
  reg [31:0] _RAND_457;
  reg [31:0] _RAND_458;
  reg [31:0] _RAND_459;
  reg [31:0] _RAND_460;
  reg [31:0] _RAND_461;
  reg [31:0] _RAND_462;
  reg [31:0] _RAND_463;
  reg [31:0] _RAND_464;
  reg [31:0] _RAND_465;
  reg [31:0] _RAND_466;
  reg [31:0] _RAND_467;
  reg [31:0] _RAND_468;
  reg [31:0] _RAND_469;
  reg [31:0] _RAND_470;
  reg [31:0] _RAND_471;
  reg [31:0] _RAND_472;
  reg [31:0] _RAND_473;
  reg [31:0] _RAND_474;
  reg [31:0] _RAND_475;
  reg [31:0] _RAND_476;
  reg [31:0] _RAND_477;
  reg [31:0] _RAND_478;
  reg [31:0] _RAND_479;
  reg [31:0] _RAND_480;
  reg [31:0] _RAND_481;
  reg [31:0] _RAND_482;
  reg [31:0] _RAND_483;
  reg [31:0] _RAND_484;
  reg [31:0] _RAND_485;
  reg [31:0] _RAND_486;
  reg [31:0] _RAND_487;
  reg [31:0] _RAND_488;
  reg [31:0] _RAND_489;
  reg [31:0] _RAND_490;
  reg [31:0] _RAND_491;
  reg [31:0] _RAND_492;
  reg [31:0] _RAND_493;
  reg [31:0] _RAND_494;
  reg [31:0] _RAND_495;
  reg [31:0] _RAND_496;
  reg [31:0] _RAND_497;
  reg [31:0] _RAND_498;
  reg [31:0] _RAND_499;
  reg [31:0] _RAND_500;
  reg [31:0] _RAND_501;
  reg [31:0] _RAND_502;
  reg [31:0] _RAND_503;
  reg [31:0] _RAND_504;
  reg [31:0] _RAND_505;
  reg [31:0] _RAND_506;
  reg [31:0] _RAND_507;
  reg [31:0] _RAND_508;
  reg [31:0] _RAND_509;
  reg [31:0] _RAND_510;
  reg [31:0] _RAND_511;
  reg [31:0] _RAND_512;
  reg [31:0] _RAND_513;
  reg [31:0] _RAND_514;
  reg [31:0] _RAND_515;
  reg [31:0] _RAND_516;
  reg [31:0] _RAND_517;
  reg [31:0] _RAND_518;
  reg [31:0] _RAND_519;
  reg [31:0] _RAND_520;
  reg [31:0] _RAND_521;
  reg [31:0] _RAND_522;
  reg [31:0] _RAND_523;
  reg [31:0] _RAND_524;
  reg [31:0] _RAND_525;
  reg [31:0] _RAND_526;
  reg [31:0] _RAND_527;
  reg [31:0] _RAND_528;
  reg [31:0] _RAND_529;
  reg [31:0] _RAND_530;
  reg [31:0] _RAND_531;
  reg [31:0] _RAND_532;
  reg [31:0] _RAND_533;
  reg [31:0] _RAND_534;
  reg [31:0] _RAND_535;
  reg [31:0] _RAND_536;
  reg [31:0] _RAND_537;
  reg [31:0] _RAND_538;
  reg [31:0] _RAND_539;
  reg [31:0] _RAND_540;
  reg [31:0] _RAND_541;
  reg [31:0] _RAND_542;
  reg [31:0] _RAND_543;
  reg [31:0] _RAND_544;
  reg [31:0] _RAND_545;
  reg [31:0] _RAND_546;
  reg [31:0] _RAND_547;
  reg [31:0] _RAND_548;
  reg [31:0] _RAND_549;
  reg [31:0] _RAND_550;
  reg [31:0] _RAND_551;
  reg [31:0] _RAND_552;
  reg [31:0] _RAND_553;
  reg [31:0] _RAND_554;
  reg [31:0] _RAND_555;
  reg [31:0] _RAND_556;
  reg [31:0] _RAND_557;
  reg [31:0] _RAND_558;
  reg [31:0] _RAND_559;
  reg [31:0] _RAND_560;
  reg [31:0] _RAND_561;
  reg [31:0] _RAND_562;
  reg [31:0] _RAND_563;
  reg [31:0] _RAND_564;
  reg [31:0] _RAND_565;
  reg [31:0] _RAND_566;
  reg [31:0] _RAND_567;
  reg [31:0] _RAND_568;
  reg [31:0] _RAND_569;
  reg [31:0] _RAND_570;
  reg [31:0] _RAND_571;
  reg [31:0] _RAND_572;
  reg [31:0] _RAND_573;
  reg [31:0] _RAND_574;
  reg [31:0] _RAND_575;
  reg [31:0] _RAND_576;
  reg [31:0] _RAND_577;
  reg [31:0] _RAND_578;
  reg [31:0] _RAND_579;
  reg [31:0] _RAND_580;
  reg [31:0] _RAND_581;
  reg [31:0] _RAND_582;
  reg [31:0] _RAND_583;
  reg [31:0] _RAND_584;
  reg [31:0] _RAND_585;
  reg [31:0] _RAND_586;
  reg [31:0] _RAND_587;
  reg [31:0] _RAND_588;
  reg [31:0] _RAND_589;
  reg [31:0] _RAND_590;
  reg [31:0] _RAND_591;
  reg [31:0] _RAND_592;
  reg [31:0] _RAND_593;
  reg [31:0] _RAND_594;
  reg [31:0] _RAND_595;
  reg [31:0] _RAND_596;
  reg [31:0] _RAND_597;
  reg [31:0] _RAND_598;
  reg [31:0] _RAND_599;
  reg [31:0] _RAND_600;
  reg [31:0] _RAND_601;
  reg [31:0] _RAND_602;
  reg [31:0] _RAND_603;
  reg [31:0] _RAND_604;
  reg [31:0] _RAND_605;
  reg [31:0] _RAND_606;
  reg [31:0] _RAND_607;
  reg [31:0] _RAND_608;
  reg [31:0] _RAND_609;
  reg [31:0] _RAND_610;
  reg [31:0] _RAND_611;
  reg [31:0] _RAND_612;
  reg [31:0] _RAND_613;
  reg [31:0] _RAND_614;
  reg [31:0] _RAND_615;
  reg [31:0] _RAND_616;
  reg [31:0] _RAND_617;
  reg [31:0] _RAND_618;
  reg [31:0] _RAND_619;
  reg [31:0] _RAND_620;
  reg [31:0] _RAND_621;
  reg [31:0] _RAND_622;
  reg [31:0] _RAND_623;
  reg [31:0] _RAND_624;
  reg [31:0] _RAND_625;
  reg [31:0] _RAND_626;
  reg [31:0] _RAND_627;
  reg [31:0] _RAND_628;
  reg [31:0] _RAND_629;
  reg [31:0] _RAND_630;
  reg [31:0] _RAND_631;
  reg [31:0] _RAND_632;
  reg [31:0] _RAND_633;
  reg [31:0] _RAND_634;
  reg [31:0] _RAND_635;
  reg [31:0] _RAND_636;
  reg [31:0] _RAND_637;
  reg [31:0] _RAND_638;
  reg [31:0] _RAND_639;
  reg [31:0] _RAND_640;
  reg [31:0] _RAND_641;
  reg [31:0] _RAND_642;
  reg [31:0] _RAND_643;
  reg [31:0] _RAND_644;
  reg [31:0] _RAND_645;
  reg [31:0] _RAND_646;
  reg [31:0] _RAND_647;
  reg [31:0] _RAND_648;
  reg [31:0] _RAND_649;
  reg [31:0] _RAND_650;
  reg [31:0] _RAND_651;
  reg [31:0] _RAND_652;
  reg [31:0] _RAND_653;
  reg [31:0] _RAND_654;
  reg [31:0] _RAND_655;
  reg [31:0] _RAND_656;
  reg [31:0] _RAND_657;
  reg [31:0] _RAND_658;
  reg [31:0] _RAND_659;
  reg [31:0] _RAND_660;
  reg [31:0] _RAND_661;
  reg [31:0] _RAND_662;
  reg [31:0] _RAND_663;
  reg [31:0] _RAND_664;
  reg [31:0] _RAND_665;
  reg [31:0] _RAND_666;
  reg [31:0] _RAND_667;
  reg [31:0] _RAND_668;
  reg [31:0] _RAND_669;
  reg [31:0] _RAND_670;
  reg [31:0] _RAND_671;
  reg [31:0] _RAND_672;
  reg [31:0] _RAND_673;
  reg [31:0] _RAND_674;
  reg [31:0] _RAND_675;
  reg [31:0] _RAND_676;
  reg [31:0] _RAND_677;
  reg [31:0] _RAND_678;
  reg [31:0] _RAND_679;
  reg [31:0] _RAND_680;
  reg [31:0] _RAND_681;
  reg [31:0] _RAND_682;
  reg [31:0] _RAND_683;
  reg [31:0] _RAND_684;
  reg [31:0] _RAND_685;
  reg [31:0] _RAND_686;
  reg [31:0] _RAND_687;
  reg [31:0] _RAND_688;
  reg [31:0] _RAND_689;
  reg [31:0] _RAND_690;
  reg [31:0] _RAND_691;
  reg [31:0] _RAND_692;
  reg [31:0] _RAND_693;
  reg [31:0] _RAND_694;
  reg [31:0] _RAND_695;
  reg [31:0] _RAND_696;
  reg [31:0] _RAND_697;
  reg [31:0] _RAND_698;
  reg [31:0] _RAND_699;
  reg [31:0] _RAND_700;
  reg [31:0] _RAND_701;
  reg [31:0] _RAND_702;
  reg [31:0] _RAND_703;
  reg [31:0] _RAND_704;
  reg [31:0] _RAND_705;
  reg [31:0] _RAND_706;
  reg [31:0] _RAND_707;
  reg [31:0] _RAND_708;
  reg [31:0] _RAND_709;
  reg [31:0] _RAND_710;
  reg [31:0] _RAND_711;
  reg [31:0] _RAND_712;
  reg [31:0] _RAND_713;
  reg [31:0] _RAND_714;
  reg [31:0] _RAND_715;
  reg [31:0] _RAND_716;
  reg [31:0] _RAND_717;
  reg [31:0] _RAND_718;
  reg [31:0] _RAND_719;
  reg [31:0] _RAND_720;
  reg [31:0] _RAND_721;
  reg [31:0] _RAND_722;
  reg [31:0] _RAND_723;
  reg [31:0] _RAND_724;
  reg [31:0] _RAND_725;
  reg [31:0] _RAND_726;
  reg [31:0] _RAND_727;
  reg [31:0] _RAND_728;
  reg [31:0] _RAND_729;
  reg [31:0] _RAND_730;
  reg [31:0] _RAND_731;
  reg [31:0] _RAND_732;
  reg [31:0] _RAND_733;
  reg [31:0] _RAND_734;
  reg [31:0] _RAND_735;
  reg [31:0] _RAND_736;
  reg [31:0] _RAND_737;
  reg [31:0] _RAND_738;
  reg [31:0] _RAND_739;
  reg [31:0] _RAND_740;
  reg [31:0] _RAND_741;
  reg [31:0] _RAND_742;
  reg [31:0] _RAND_743;
  reg [31:0] _RAND_744;
  reg [31:0] _RAND_745;
  reg [31:0] _RAND_746;
  reg [31:0] _RAND_747;
  reg [31:0] _RAND_748;
  reg [31:0] _RAND_749;
  reg [31:0] _RAND_750;
  reg [31:0] _RAND_751;
  reg [31:0] _RAND_752;
  reg [31:0] _RAND_753;
  reg [31:0] _RAND_754;
  reg [31:0] _RAND_755;
  reg [31:0] _RAND_756;
  reg [31:0] _RAND_757;
  reg [31:0] _RAND_758;
  reg [31:0] _RAND_759;
  reg [31:0] _RAND_760;
  reg [31:0] _RAND_761;
  reg [31:0] _RAND_762;
  reg [31:0] _RAND_763;
  reg [31:0] _RAND_764;
  reg [31:0] _RAND_765;
  reg [31:0] _RAND_766;
  reg [31:0] _RAND_767;
  reg [31:0] _RAND_768;
  reg [31:0] _RAND_769;
  reg [31:0] _RAND_770;
  reg [31:0] _RAND_771;
  reg [31:0] _RAND_772;
  reg [31:0] _RAND_773;
  reg [31:0] _RAND_774;
  reg [31:0] _RAND_775;
  reg [31:0] _RAND_776;
  reg [31:0] _RAND_777;
  reg [31:0] _RAND_778;
  reg [31:0] _RAND_779;
  reg [31:0] _RAND_780;
  reg [31:0] _RAND_781;
  reg [31:0] _RAND_782;
  reg [31:0] _RAND_783;
`endif // RANDOMIZE_REG_INIT
  wire [7:0] MulAdd_io__b_0; // @[ChiselImProc.scala 244:29]
  wire [7:0] MulAdd_io__b_1; // @[ChiselImProc.scala 244:29]
  wire [7:0] MulAdd_io__b_2; // @[ChiselImProc.scala 244:29]
  wire [7:0] MulAdd_io__b_3; // @[ChiselImProc.scala 244:29]
  wire [7:0] MulAdd_io__b_4; // @[ChiselImProc.scala 244:29]
  wire [7:0] MulAdd_io__b_5; // @[ChiselImProc.scala 244:29]
  wire [7:0] MulAdd_io__b_6; // @[ChiselImProc.scala 244:29]
  wire [7:0] MulAdd_io__b_7; // @[ChiselImProc.scala 244:29]
  wire [7:0] MulAdd_io__b_8; // @[ChiselImProc.scala 244:29]
  wire [15:0] MulAdd_io__output; // @[ChiselImProc.scala 244:29]
  wire [15:0] MulAdd_io_output; // @[ChiselImProc.scala 244:29]
  reg [1:0] stateReg; // @[ChiselImProc.scala 62:28]
  reg [7:0] dataReg; // @[ChiselImProc.scala 64:23]
  reg [7:0] shadowReg; // @[ChiselImProc.scala 66:25]
  reg  userReg; // @[ChiselImProc.scala 67:23]
  reg  shadowUserReg; // @[ChiselImProc.scala 68:29]
  reg  lastReg; // @[ChiselImProc.scala 69:23]
  reg  shadowLastReg; // @[ChiselImProc.scala 70:29]
  wire  _T = 2'h0 == stateReg; // @[Conditional.scala 37:30]
  wire  _T_1 = 2'h1 == stateReg; // @[Conditional.scala 37:30]
  wire  _T_2 = ~io__enq_valid; // @[ChiselImProc.scala 84:39]
  wire  _T_3 = io__deq_ready & _T_2; // @[ChiselImProc.scala 84:36]
  wire  _T_4 = io__deq_ready & io__enq_valid; // @[ChiselImProc.scala 87:42]
  wire  _T_5 = ~io__deq_ready; // @[ChiselImProc.scala 92:29]
  wire  _T_6 = _T_5 & io__enq_valid; // @[ChiselImProc.scala 92:43]
  wire  _T_7 = 2'h2 == stateReg; // @[Conditional.scala 37:30]
  wire  _T_8 = 2'h3 == stateReg; // @[Conditional.scala 37:30]
  wire  _T_9 = stateReg == 2'h0; // @[ChiselImProc.scala 116:35]
  wire  _T_10 = stateReg == 2'h1; // @[ChiselImProc.scala 116:57]
  wire  _T_11 = _T_9 | _T_10; // @[ChiselImProc.scala 116:45]
  wire  _T_12 = stateReg == 2'h3; // @[ChiselImProc.scala 116:77]
  wire  _T_15 = stateReg == 2'h2; // @[ChiselImProc.scala 117:55]
  wire  _T_16 = _T_10 | _T_15; // @[ChiselImProc.scala 117:43]
  reg [7:0] lineBuffer_0; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_1; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_2; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_3; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_4; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_5; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_6; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_7; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_8; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_9; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_10; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_11; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_12; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_13; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_14; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_15; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_16; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_17; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_18; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_19; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_20; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_21; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_22; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_23; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_24; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_25; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_26; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_27; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_28; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_29; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_30; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_31; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_32; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_33; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_34; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_35; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_36; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_37; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_38; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_39; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_40; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_41; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_42; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_43; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_44; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_45; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_46; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_47; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_48; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_49; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_50; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_51; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_52; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_53; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_54; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_55; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_56; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_57; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_58; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_59; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_60; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_61; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_62; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_63; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_64; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_65; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_66; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_67; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_68; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_69; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_70; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_71; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_72; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_73; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_74; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_75; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_76; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_77; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_78; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_79; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_80; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_81; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_82; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_83; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_84; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_85; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_86; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_87; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_88; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_89; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_90; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_91; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_92; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_93; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_94; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_95; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_96; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_97; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_98; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_99; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_100; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_101; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_102; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_103; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_104; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_105; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_106; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_107; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_108; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_109; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_110; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_111; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_112; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_113; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_114; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_115; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_116; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_117; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_118; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_119; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_120; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_121; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_122; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_123; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_124; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_125; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_126; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_127; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_128; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_129; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_130; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_131; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_132; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_133; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_134; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_135; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_136; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_137; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_138; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_139; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_140; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_141; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_142; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_143; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_144; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_145; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_146; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_147; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_148; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_149; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_150; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_151; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_152; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_153; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_154; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_155; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_156; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_157; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_158; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_159; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_160; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_161; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_162; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_163; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_164; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_165; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_166; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_167; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_168; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_169; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_170; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_171; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_172; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_173; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_174; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_175; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_176; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_177; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_178; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_179; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_180; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_181; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_182; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_183; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_184; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_185; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_186; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_187; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_188; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_189; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_190; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_191; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_192; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_193; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_194; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_195; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_196; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_197; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_198; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_199; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_200; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_201; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_202; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_203; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_204; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_205; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_206; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_207; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_208; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_209; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_210; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_211; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_212; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_213; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_214; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_215; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_216; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_217; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_218; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_219; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_220; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_221; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_222; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_223; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_224; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_225; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_226; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_227; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_228; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_229; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_230; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_231; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_232; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_233; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_234; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_235; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_236; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_237; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_238; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_239; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_240; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_241; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_242; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_243; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_244; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_245; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_246; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_247; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_248; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_249; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_250; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_251; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_252; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_253; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_254; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_255; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_256; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_257; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_258; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_259; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_260; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_261; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_262; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_263; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_264; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_265; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_266; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_267; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_268; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_269; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_270; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_271; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_272; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_273; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_274; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_275; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_276; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_277; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_278; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_279; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_280; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_281; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_282; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_283; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_284; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_285; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_286; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_287; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_288; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_289; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_290; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_291; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_292; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_293; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_294; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_295; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_296; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_297; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_298; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_299; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_300; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_301; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_302; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_303; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_304; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_305; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_306; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_307; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_308; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_309; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_310; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_311; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_312; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_313; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_314; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_315; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_316; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_317; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_318; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_319; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_320; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_321; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_322; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_323; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_324; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_325; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_326; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_327; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_328; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_329; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_330; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_331; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_332; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_333; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_334; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_335; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_336; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_337; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_338; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_339; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_340; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_341; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_342; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_343; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_344; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_345; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_346; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_347; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_348; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_349; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_350; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_351; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_352; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_353; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_354; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_355; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_356; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_357; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_358; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_359; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_360; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_361; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_362; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_363; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_364; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_365; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_366; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_367; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_368; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_369; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_370; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_371; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_372; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_373; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_374; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_375; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_376; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_377; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_378; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_379; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_380; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_381; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_382; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_383; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_384; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_385; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_386; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_387; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_388; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_389; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_390; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_391; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_392; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_393; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_394; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_395; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_396; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_397; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_398; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_399; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_400; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_401; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_402; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_403; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_404; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_405; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_406; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_407; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_408; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_409; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_410; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_411; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_412; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_413; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_414; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_415; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_416; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_417; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_418; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_419; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_420; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_421; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_422; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_423; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_424; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_425; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_426; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_427; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_428; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_429; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_430; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_431; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_432; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_433; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_434; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_435; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_436; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_437; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_438; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_439; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_440; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_441; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_442; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_443; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_444; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_445; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_446; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_447; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_448; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_449; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_450; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_451; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_452; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_453; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_454; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_455; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_456; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_457; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_458; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_459; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_460; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_461; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_462; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_463; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_464; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_465; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_466; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_467; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_468; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_469; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_470; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_471; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_472; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_473; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_474; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_475; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_476; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_477; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_478; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_479; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_480; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_481; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_482; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_483; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_484; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_485; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_486; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_487; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_488; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_489; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_490; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_491; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_492; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_493; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_494; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_495; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_496; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_497; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_498; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_499; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_500; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_501; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_502; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_503; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_504; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_505; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_506; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_507; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_508; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_509; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_510; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_511; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_512; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_513; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_514; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_515; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_516; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_517; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_518; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_519; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_520; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_521; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_522; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_523; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_524; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_525; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_526; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_527; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_528; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_529; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_530; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_531; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_532; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_533; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_534; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_535; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_536; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_537; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_538; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_539; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_540; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_541; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_542; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_543; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_544; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_545; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_546; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_547; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_548; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_549; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_550; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_551; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_552; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_553; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_554; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_555; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_556; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_557; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_558; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_559; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_560; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_561; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_562; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_563; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_564; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_565; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_566; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_567; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_568; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_569; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_570; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_571; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_572; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_573; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_574; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_575; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_576; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_577; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_578; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_579; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_580; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_581; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_582; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_583; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_584; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_585; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_586; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_587; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_588; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_589; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_590; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_591; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_592; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_593; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_594; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_595; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_596; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_597; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_598; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_599; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_600; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_601; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_602; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_603; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_604; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_605; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_606; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_607; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_608; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_609; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_610; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_611; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_612; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_613; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_614; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_615; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_616; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_617; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_618; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_619; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_620; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_621; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_622; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_623; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_624; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_625; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_626; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_627; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_628; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_629; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_630; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_631; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_632; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_633; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_634; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_635; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_636; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_637; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_638; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_639; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_640; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_641; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_642; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_643; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_644; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_645; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_646; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_647; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_648; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_649; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_650; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_651; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_652; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_653; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_654; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_655; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_656; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_657; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_658; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_659; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_660; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_661; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_662; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_663; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_664; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_665; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_666; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_667; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_668; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_669; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_670; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_671; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_672; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_673; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_674; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_675; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_676; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_677; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_678; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_679; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_680; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_681; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_682; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_683; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_684; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_685; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_686; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_687; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_688; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_689; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_690; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_691; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_692; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_693; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_694; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_695; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_696; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_697; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_698; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_699; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_700; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_701; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_702; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_703; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_704; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_705; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_706; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_707; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_708; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_709; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_710; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_711; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_712; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_713; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_714; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_715; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_716; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_717; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_718; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_719; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_720; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_721; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_722; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_723; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_724; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_725; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_726; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_727; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_728; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_729; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_730; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_731; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_732; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_733; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_734; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_735; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_736; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_737; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_738; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_739; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_740; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_741; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_742; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_743; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_744; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_745; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_746; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_747; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_748; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_749; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_750; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_751; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_752; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_753; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_754; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_755; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_756; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_757; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_758; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_759; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_760; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_761; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_762; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_763; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_764; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_765; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_766; // @[ChiselImProc.scala 226:26]
  reg [7:0] lineBuffer_767; // @[ChiselImProc.scala 226:26]
  reg [7:0] windowBuffer_0; // @[ChiselImProc.scala 227:28]
  reg [7:0] windowBuffer_1; // @[ChiselImProc.scala 227:28]
  reg [7:0] windowBuffer_2; // @[ChiselImProc.scala 227:28]
  reg [7:0] windowBuffer_3; // @[ChiselImProc.scala 227:28]
  reg [7:0] windowBuffer_4; // @[ChiselImProc.scala 227:28]
  reg [7:0] windowBuffer_5; // @[ChiselImProc.scala 227:28]
  reg [7:0] windowBuffer_6; // @[ChiselImProc.scala 227:28]
  reg [7:0] windowBuffer_7; // @[ChiselImProc.scala 227:28]
  reg [7:0] windowBuffer_8; // @[ChiselImProc.scala 227:28]
  wire  sel = _T_16 & io__deq_ready; // @[ChiselImProc.scala 230:47]
  wire [71:0] _T_805 = {windowBuffer_0,windowBuffer_1,windowBuffer_2,windowBuffer_3,windowBuffer_4,windowBuffer_5,windowBuffer_6,windowBuffer_7,windowBuffer_8}; // @[Cat.scala 29:58]
  MulAdd MulAdd ( // @[ChiselImProc.scala 244:29]
    .io__b_0(MulAdd_io__b_0),
    .io__b_1(MulAdd_io__b_1),
    .io__b_2(MulAdd_io__b_2),
    .io__b_3(MulAdd_io__b_3),
    .io__b_4(MulAdd_io__b_4),
    .io__b_5(MulAdd_io__b_5),
    .io__b_6(MulAdd_io__b_6),
    .io__b_7(MulAdd_io__b_7),
    .io__b_8(MulAdd_io__b_8),
    .io__output(MulAdd_io__output),
    .io_output(MulAdd_io_output)
  );
  assign io__enq_ready = _T_11 | _T_12; // @[ChiselImProc.scala 116:22]
  assign io__deq_valid = _T_10 | _T_15; // @[ChiselImProc.scala 117:22]
  assign io__deq_bits = MulAdd_io__output[11:4]; // @[ChiselImProc.scala 254:17]
  assign io__deq_user = userReg; // @[ChiselImProc.scala 144:17 ChiselImProc.scala 114:21]
  assign io__deq_last = lastReg; // @[ChiselImProc.scala 143:17 ChiselImProc.scala 113:21]
  assign io_deq_ready = io__deq_ready;
  assign io_deq_valid = io__deq_valid;
  assign _T_805_0 = _T_805;
  assign io_output = MulAdd_io_output;
  assign MulAdd_io__b_0 = windowBuffer_0; // @[ChiselImProc.scala 252:13]
  assign MulAdd_io__b_1 = windowBuffer_1; // @[ChiselImProc.scala 252:13]
  assign MulAdd_io__b_2 = windowBuffer_2; // @[ChiselImProc.scala 252:13]
  assign MulAdd_io__b_3 = windowBuffer_3; // @[ChiselImProc.scala 252:13]
  assign MulAdd_io__b_4 = windowBuffer_4; // @[ChiselImProc.scala 252:13]
  assign MulAdd_io__b_5 = windowBuffer_5; // @[ChiselImProc.scala 252:13]
  assign MulAdd_io__b_6 = windowBuffer_6; // @[ChiselImProc.scala 252:13]
  assign MulAdd_io__b_7 = windowBuffer_7; // @[ChiselImProc.scala 252:13]
  assign MulAdd_io__b_8 = windowBuffer_8; // @[ChiselImProc.scala 252:13]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  stateReg = _RAND_0[1:0];
  _RAND_1 = {1{`RANDOM}};
  dataReg = _RAND_1[7:0];
  _RAND_2 = {1{`RANDOM}};
  shadowReg = _RAND_2[7:0];
  _RAND_3 = {1{`RANDOM}};
  userReg = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  shadowUserReg = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  lastReg = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  shadowLastReg = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  lineBuffer_0 = _RAND_7[7:0];
  _RAND_8 = {1{`RANDOM}};
  lineBuffer_1 = _RAND_8[7:0];
  _RAND_9 = {1{`RANDOM}};
  lineBuffer_2 = _RAND_9[7:0];
  _RAND_10 = {1{`RANDOM}};
  lineBuffer_3 = _RAND_10[7:0];
  _RAND_11 = {1{`RANDOM}};
  lineBuffer_4 = _RAND_11[7:0];
  _RAND_12 = {1{`RANDOM}};
  lineBuffer_5 = _RAND_12[7:0];
  _RAND_13 = {1{`RANDOM}};
  lineBuffer_6 = _RAND_13[7:0];
  _RAND_14 = {1{`RANDOM}};
  lineBuffer_7 = _RAND_14[7:0];
  _RAND_15 = {1{`RANDOM}};
  lineBuffer_8 = _RAND_15[7:0];
  _RAND_16 = {1{`RANDOM}};
  lineBuffer_9 = _RAND_16[7:0];
  _RAND_17 = {1{`RANDOM}};
  lineBuffer_10 = _RAND_17[7:0];
  _RAND_18 = {1{`RANDOM}};
  lineBuffer_11 = _RAND_18[7:0];
  _RAND_19 = {1{`RANDOM}};
  lineBuffer_12 = _RAND_19[7:0];
  _RAND_20 = {1{`RANDOM}};
  lineBuffer_13 = _RAND_20[7:0];
  _RAND_21 = {1{`RANDOM}};
  lineBuffer_14 = _RAND_21[7:0];
  _RAND_22 = {1{`RANDOM}};
  lineBuffer_15 = _RAND_22[7:0];
  _RAND_23 = {1{`RANDOM}};
  lineBuffer_16 = _RAND_23[7:0];
  _RAND_24 = {1{`RANDOM}};
  lineBuffer_17 = _RAND_24[7:0];
  _RAND_25 = {1{`RANDOM}};
  lineBuffer_18 = _RAND_25[7:0];
  _RAND_26 = {1{`RANDOM}};
  lineBuffer_19 = _RAND_26[7:0];
  _RAND_27 = {1{`RANDOM}};
  lineBuffer_20 = _RAND_27[7:0];
  _RAND_28 = {1{`RANDOM}};
  lineBuffer_21 = _RAND_28[7:0];
  _RAND_29 = {1{`RANDOM}};
  lineBuffer_22 = _RAND_29[7:0];
  _RAND_30 = {1{`RANDOM}};
  lineBuffer_23 = _RAND_30[7:0];
  _RAND_31 = {1{`RANDOM}};
  lineBuffer_24 = _RAND_31[7:0];
  _RAND_32 = {1{`RANDOM}};
  lineBuffer_25 = _RAND_32[7:0];
  _RAND_33 = {1{`RANDOM}};
  lineBuffer_26 = _RAND_33[7:0];
  _RAND_34 = {1{`RANDOM}};
  lineBuffer_27 = _RAND_34[7:0];
  _RAND_35 = {1{`RANDOM}};
  lineBuffer_28 = _RAND_35[7:0];
  _RAND_36 = {1{`RANDOM}};
  lineBuffer_29 = _RAND_36[7:0];
  _RAND_37 = {1{`RANDOM}};
  lineBuffer_30 = _RAND_37[7:0];
  _RAND_38 = {1{`RANDOM}};
  lineBuffer_31 = _RAND_38[7:0];
  _RAND_39 = {1{`RANDOM}};
  lineBuffer_32 = _RAND_39[7:0];
  _RAND_40 = {1{`RANDOM}};
  lineBuffer_33 = _RAND_40[7:0];
  _RAND_41 = {1{`RANDOM}};
  lineBuffer_34 = _RAND_41[7:0];
  _RAND_42 = {1{`RANDOM}};
  lineBuffer_35 = _RAND_42[7:0];
  _RAND_43 = {1{`RANDOM}};
  lineBuffer_36 = _RAND_43[7:0];
  _RAND_44 = {1{`RANDOM}};
  lineBuffer_37 = _RAND_44[7:0];
  _RAND_45 = {1{`RANDOM}};
  lineBuffer_38 = _RAND_45[7:0];
  _RAND_46 = {1{`RANDOM}};
  lineBuffer_39 = _RAND_46[7:0];
  _RAND_47 = {1{`RANDOM}};
  lineBuffer_40 = _RAND_47[7:0];
  _RAND_48 = {1{`RANDOM}};
  lineBuffer_41 = _RAND_48[7:0];
  _RAND_49 = {1{`RANDOM}};
  lineBuffer_42 = _RAND_49[7:0];
  _RAND_50 = {1{`RANDOM}};
  lineBuffer_43 = _RAND_50[7:0];
  _RAND_51 = {1{`RANDOM}};
  lineBuffer_44 = _RAND_51[7:0];
  _RAND_52 = {1{`RANDOM}};
  lineBuffer_45 = _RAND_52[7:0];
  _RAND_53 = {1{`RANDOM}};
  lineBuffer_46 = _RAND_53[7:0];
  _RAND_54 = {1{`RANDOM}};
  lineBuffer_47 = _RAND_54[7:0];
  _RAND_55 = {1{`RANDOM}};
  lineBuffer_48 = _RAND_55[7:0];
  _RAND_56 = {1{`RANDOM}};
  lineBuffer_49 = _RAND_56[7:0];
  _RAND_57 = {1{`RANDOM}};
  lineBuffer_50 = _RAND_57[7:0];
  _RAND_58 = {1{`RANDOM}};
  lineBuffer_51 = _RAND_58[7:0];
  _RAND_59 = {1{`RANDOM}};
  lineBuffer_52 = _RAND_59[7:0];
  _RAND_60 = {1{`RANDOM}};
  lineBuffer_53 = _RAND_60[7:0];
  _RAND_61 = {1{`RANDOM}};
  lineBuffer_54 = _RAND_61[7:0];
  _RAND_62 = {1{`RANDOM}};
  lineBuffer_55 = _RAND_62[7:0];
  _RAND_63 = {1{`RANDOM}};
  lineBuffer_56 = _RAND_63[7:0];
  _RAND_64 = {1{`RANDOM}};
  lineBuffer_57 = _RAND_64[7:0];
  _RAND_65 = {1{`RANDOM}};
  lineBuffer_58 = _RAND_65[7:0];
  _RAND_66 = {1{`RANDOM}};
  lineBuffer_59 = _RAND_66[7:0];
  _RAND_67 = {1{`RANDOM}};
  lineBuffer_60 = _RAND_67[7:0];
  _RAND_68 = {1{`RANDOM}};
  lineBuffer_61 = _RAND_68[7:0];
  _RAND_69 = {1{`RANDOM}};
  lineBuffer_62 = _RAND_69[7:0];
  _RAND_70 = {1{`RANDOM}};
  lineBuffer_63 = _RAND_70[7:0];
  _RAND_71 = {1{`RANDOM}};
  lineBuffer_64 = _RAND_71[7:0];
  _RAND_72 = {1{`RANDOM}};
  lineBuffer_65 = _RAND_72[7:0];
  _RAND_73 = {1{`RANDOM}};
  lineBuffer_66 = _RAND_73[7:0];
  _RAND_74 = {1{`RANDOM}};
  lineBuffer_67 = _RAND_74[7:0];
  _RAND_75 = {1{`RANDOM}};
  lineBuffer_68 = _RAND_75[7:0];
  _RAND_76 = {1{`RANDOM}};
  lineBuffer_69 = _RAND_76[7:0];
  _RAND_77 = {1{`RANDOM}};
  lineBuffer_70 = _RAND_77[7:0];
  _RAND_78 = {1{`RANDOM}};
  lineBuffer_71 = _RAND_78[7:0];
  _RAND_79 = {1{`RANDOM}};
  lineBuffer_72 = _RAND_79[7:0];
  _RAND_80 = {1{`RANDOM}};
  lineBuffer_73 = _RAND_80[7:0];
  _RAND_81 = {1{`RANDOM}};
  lineBuffer_74 = _RAND_81[7:0];
  _RAND_82 = {1{`RANDOM}};
  lineBuffer_75 = _RAND_82[7:0];
  _RAND_83 = {1{`RANDOM}};
  lineBuffer_76 = _RAND_83[7:0];
  _RAND_84 = {1{`RANDOM}};
  lineBuffer_77 = _RAND_84[7:0];
  _RAND_85 = {1{`RANDOM}};
  lineBuffer_78 = _RAND_85[7:0];
  _RAND_86 = {1{`RANDOM}};
  lineBuffer_79 = _RAND_86[7:0];
  _RAND_87 = {1{`RANDOM}};
  lineBuffer_80 = _RAND_87[7:0];
  _RAND_88 = {1{`RANDOM}};
  lineBuffer_81 = _RAND_88[7:0];
  _RAND_89 = {1{`RANDOM}};
  lineBuffer_82 = _RAND_89[7:0];
  _RAND_90 = {1{`RANDOM}};
  lineBuffer_83 = _RAND_90[7:0];
  _RAND_91 = {1{`RANDOM}};
  lineBuffer_84 = _RAND_91[7:0];
  _RAND_92 = {1{`RANDOM}};
  lineBuffer_85 = _RAND_92[7:0];
  _RAND_93 = {1{`RANDOM}};
  lineBuffer_86 = _RAND_93[7:0];
  _RAND_94 = {1{`RANDOM}};
  lineBuffer_87 = _RAND_94[7:0];
  _RAND_95 = {1{`RANDOM}};
  lineBuffer_88 = _RAND_95[7:0];
  _RAND_96 = {1{`RANDOM}};
  lineBuffer_89 = _RAND_96[7:0];
  _RAND_97 = {1{`RANDOM}};
  lineBuffer_90 = _RAND_97[7:0];
  _RAND_98 = {1{`RANDOM}};
  lineBuffer_91 = _RAND_98[7:0];
  _RAND_99 = {1{`RANDOM}};
  lineBuffer_92 = _RAND_99[7:0];
  _RAND_100 = {1{`RANDOM}};
  lineBuffer_93 = _RAND_100[7:0];
  _RAND_101 = {1{`RANDOM}};
  lineBuffer_94 = _RAND_101[7:0];
  _RAND_102 = {1{`RANDOM}};
  lineBuffer_95 = _RAND_102[7:0];
  _RAND_103 = {1{`RANDOM}};
  lineBuffer_96 = _RAND_103[7:0];
  _RAND_104 = {1{`RANDOM}};
  lineBuffer_97 = _RAND_104[7:0];
  _RAND_105 = {1{`RANDOM}};
  lineBuffer_98 = _RAND_105[7:0];
  _RAND_106 = {1{`RANDOM}};
  lineBuffer_99 = _RAND_106[7:0];
  _RAND_107 = {1{`RANDOM}};
  lineBuffer_100 = _RAND_107[7:0];
  _RAND_108 = {1{`RANDOM}};
  lineBuffer_101 = _RAND_108[7:0];
  _RAND_109 = {1{`RANDOM}};
  lineBuffer_102 = _RAND_109[7:0];
  _RAND_110 = {1{`RANDOM}};
  lineBuffer_103 = _RAND_110[7:0];
  _RAND_111 = {1{`RANDOM}};
  lineBuffer_104 = _RAND_111[7:0];
  _RAND_112 = {1{`RANDOM}};
  lineBuffer_105 = _RAND_112[7:0];
  _RAND_113 = {1{`RANDOM}};
  lineBuffer_106 = _RAND_113[7:0];
  _RAND_114 = {1{`RANDOM}};
  lineBuffer_107 = _RAND_114[7:0];
  _RAND_115 = {1{`RANDOM}};
  lineBuffer_108 = _RAND_115[7:0];
  _RAND_116 = {1{`RANDOM}};
  lineBuffer_109 = _RAND_116[7:0];
  _RAND_117 = {1{`RANDOM}};
  lineBuffer_110 = _RAND_117[7:0];
  _RAND_118 = {1{`RANDOM}};
  lineBuffer_111 = _RAND_118[7:0];
  _RAND_119 = {1{`RANDOM}};
  lineBuffer_112 = _RAND_119[7:0];
  _RAND_120 = {1{`RANDOM}};
  lineBuffer_113 = _RAND_120[7:0];
  _RAND_121 = {1{`RANDOM}};
  lineBuffer_114 = _RAND_121[7:0];
  _RAND_122 = {1{`RANDOM}};
  lineBuffer_115 = _RAND_122[7:0];
  _RAND_123 = {1{`RANDOM}};
  lineBuffer_116 = _RAND_123[7:0];
  _RAND_124 = {1{`RANDOM}};
  lineBuffer_117 = _RAND_124[7:0];
  _RAND_125 = {1{`RANDOM}};
  lineBuffer_118 = _RAND_125[7:0];
  _RAND_126 = {1{`RANDOM}};
  lineBuffer_119 = _RAND_126[7:0];
  _RAND_127 = {1{`RANDOM}};
  lineBuffer_120 = _RAND_127[7:0];
  _RAND_128 = {1{`RANDOM}};
  lineBuffer_121 = _RAND_128[7:0];
  _RAND_129 = {1{`RANDOM}};
  lineBuffer_122 = _RAND_129[7:0];
  _RAND_130 = {1{`RANDOM}};
  lineBuffer_123 = _RAND_130[7:0];
  _RAND_131 = {1{`RANDOM}};
  lineBuffer_124 = _RAND_131[7:0];
  _RAND_132 = {1{`RANDOM}};
  lineBuffer_125 = _RAND_132[7:0];
  _RAND_133 = {1{`RANDOM}};
  lineBuffer_126 = _RAND_133[7:0];
  _RAND_134 = {1{`RANDOM}};
  lineBuffer_127 = _RAND_134[7:0];
  _RAND_135 = {1{`RANDOM}};
  lineBuffer_128 = _RAND_135[7:0];
  _RAND_136 = {1{`RANDOM}};
  lineBuffer_129 = _RAND_136[7:0];
  _RAND_137 = {1{`RANDOM}};
  lineBuffer_130 = _RAND_137[7:0];
  _RAND_138 = {1{`RANDOM}};
  lineBuffer_131 = _RAND_138[7:0];
  _RAND_139 = {1{`RANDOM}};
  lineBuffer_132 = _RAND_139[7:0];
  _RAND_140 = {1{`RANDOM}};
  lineBuffer_133 = _RAND_140[7:0];
  _RAND_141 = {1{`RANDOM}};
  lineBuffer_134 = _RAND_141[7:0];
  _RAND_142 = {1{`RANDOM}};
  lineBuffer_135 = _RAND_142[7:0];
  _RAND_143 = {1{`RANDOM}};
  lineBuffer_136 = _RAND_143[7:0];
  _RAND_144 = {1{`RANDOM}};
  lineBuffer_137 = _RAND_144[7:0];
  _RAND_145 = {1{`RANDOM}};
  lineBuffer_138 = _RAND_145[7:0];
  _RAND_146 = {1{`RANDOM}};
  lineBuffer_139 = _RAND_146[7:0];
  _RAND_147 = {1{`RANDOM}};
  lineBuffer_140 = _RAND_147[7:0];
  _RAND_148 = {1{`RANDOM}};
  lineBuffer_141 = _RAND_148[7:0];
  _RAND_149 = {1{`RANDOM}};
  lineBuffer_142 = _RAND_149[7:0];
  _RAND_150 = {1{`RANDOM}};
  lineBuffer_143 = _RAND_150[7:0];
  _RAND_151 = {1{`RANDOM}};
  lineBuffer_144 = _RAND_151[7:0];
  _RAND_152 = {1{`RANDOM}};
  lineBuffer_145 = _RAND_152[7:0];
  _RAND_153 = {1{`RANDOM}};
  lineBuffer_146 = _RAND_153[7:0];
  _RAND_154 = {1{`RANDOM}};
  lineBuffer_147 = _RAND_154[7:0];
  _RAND_155 = {1{`RANDOM}};
  lineBuffer_148 = _RAND_155[7:0];
  _RAND_156 = {1{`RANDOM}};
  lineBuffer_149 = _RAND_156[7:0];
  _RAND_157 = {1{`RANDOM}};
  lineBuffer_150 = _RAND_157[7:0];
  _RAND_158 = {1{`RANDOM}};
  lineBuffer_151 = _RAND_158[7:0];
  _RAND_159 = {1{`RANDOM}};
  lineBuffer_152 = _RAND_159[7:0];
  _RAND_160 = {1{`RANDOM}};
  lineBuffer_153 = _RAND_160[7:0];
  _RAND_161 = {1{`RANDOM}};
  lineBuffer_154 = _RAND_161[7:0];
  _RAND_162 = {1{`RANDOM}};
  lineBuffer_155 = _RAND_162[7:0];
  _RAND_163 = {1{`RANDOM}};
  lineBuffer_156 = _RAND_163[7:0];
  _RAND_164 = {1{`RANDOM}};
  lineBuffer_157 = _RAND_164[7:0];
  _RAND_165 = {1{`RANDOM}};
  lineBuffer_158 = _RAND_165[7:0];
  _RAND_166 = {1{`RANDOM}};
  lineBuffer_159 = _RAND_166[7:0];
  _RAND_167 = {1{`RANDOM}};
  lineBuffer_160 = _RAND_167[7:0];
  _RAND_168 = {1{`RANDOM}};
  lineBuffer_161 = _RAND_168[7:0];
  _RAND_169 = {1{`RANDOM}};
  lineBuffer_162 = _RAND_169[7:0];
  _RAND_170 = {1{`RANDOM}};
  lineBuffer_163 = _RAND_170[7:0];
  _RAND_171 = {1{`RANDOM}};
  lineBuffer_164 = _RAND_171[7:0];
  _RAND_172 = {1{`RANDOM}};
  lineBuffer_165 = _RAND_172[7:0];
  _RAND_173 = {1{`RANDOM}};
  lineBuffer_166 = _RAND_173[7:0];
  _RAND_174 = {1{`RANDOM}};
  lineBuffer_167 = _RAND_174[7:0];
  _RAND_175 = {1{`RANDOM}};
  lineBuffer_168 = _RAND_175[7:0];
  _RAND_176 = {1{`RANDOM}};
  lineBuffer_169 = _RAND_176[7:0];
  _RAND_177 = {1{`RANDOM}};
  lineBuffer_170 = _RAND_177[7:0];
  _RAND_178 = {1{`RANDOM}};
  lineBuffer_171 = _RAND_178[7:0];
  _RAND_179 = {1{`RANDOM}};
  lineBuffer_172 = _RAND_179[7:0];
  _RAND_180 = {1{`RANDOM}};
  lineBuffer_173 = _RAND_180[7:0];
  _RAND_181 = {1{`RANDOM}};
  lineBuffer_174 = _RAND_181[7:0];
  _RAND_182 = {1{`RANDOM}};
  lineBuffer_175 = _RAND_182[7:0];
  _RAND_183 = {1{`RANDOM}};
  lineBuffer_176 = _RAND_183[7:0];
  _RAND_184 = {1{`RANDOM}};
  lineBuffer_177 = _RAND_184[7:0];
  _RAND_185 = {1{`RANDOM}};
  lineBuffer_178 = _RAND_185[7:0];
  _RAND_186 = {1{`RANDOM}};
  lineBuffer_179 = _RAND_186[7:0];
  _RAND_187 = {1{`RANDOM}};
  lineBuffer_180 = _RAND_187[7:0];
  _RAND_188 = {1{`RANDOM}};
  lineBuffer_181 = _RAND_188[7:0];
  _RAND_189 = {1{`RANDOM}};
  lineBuffer_182 = _RAND_189[7:0];
  _RAND_190 = {1{`RANDOM}};
  lineBuffer_183 = _RAND_190[7:0];
  _RAND_191 = {1{`RANDOM}};
  lineBuffer_184 = _RAND_191[7:0];
  _RAND_192 = {1{`RANDOM}};
  lineBuffer_185 = _RAND_192[7:0];
  _RAND_193 = {1{`RANDOM}};
  lineBuffer_186 = _RAND_193[7:0];
  _RAND_194 = {1{`RANDOM}};
  lineBuffer_187 = _RAND_194[7:0];
  _RAND_195 = {1{`RANDOM}};
  lineBuffer_188 = _RAND_195[7:0];
  _RAND_196 = {1{`RANDOM}};
  lineBuffer_189 = _RAND_196[7:0];
  _RAND_197 = {1{`RANDOM}};
  lineBuffer_190 = _RAND_197[7:0];
  _RAND_198 = {1{`RANDOM}};
  lineBuffer_191 = _RAND_198[7:0];
  _RAND_199 = {1{`RANDOM}};
  lineBuffer_192 = _RAND_199[7:0];
  _RAND_200 = {1{`RANDOM}};
  lineBuffer_193 = _RAND_200[7:0];
  _RAND_201 = {1{`RANDOM}};
  lineBuffer_194 = _RAND_201[7:0];
  _RAND_202 = {1{`RANDOM}};
  lineBuffer_195 = _RAND_202[7:0];
  _RAND_203 = {1{`RANDOM}};
  lineBuffer_196 = _RAND_203[7:0];
  _RAND_204 = {1{`RANDOM}};
  lineBuffer_197 = _RAND_204[7:0];
  _RAND_205 = {1{`RANDOM}};
  lineBuffer_198 = _RAND_205[7:0];
  _RAND_206 = {1{`RANDOM}};
  lineBuffer_199 = _RAND_206[7:0];
  _RAND_207 = {1{`RANDOM}};
  lineBuffer_200 = _RAND_207[7:0];
  _RAND_208 = {1{`RANDOM}};
  lineBuffer_201 = _RAND_208[7:0];
  _RAND_209 = {1{`RANDOM}};
  lineBuffer_202 = _RAND_209[7:0];
  _RAND_210 = {1{`RANDOM}};
  lineBuffer_203 = _RAND_210[7:0];
  _RAND_211 = {1{`RANDOM}};
  lineBuffer_204 = _RAND_211[7:0];
  _RAND_212 = {1{`RANDOM}};
  lineBuffer_205 = _RAND_212[7:0];
  _RAND_213 = {1{`RANDOM}};
  lineBuffer_206 = _RAND_213[7:0];
  _RAND_214 = {1{`RANDOM}};
  lineBuffer_207 = _RAND_214[7:0];
  _RAND_215 = {1{`RANDOM}};
  lineBuffer_208 = _RAND_215[7:0];
  _RAND_216 = {1{`RANDOM}};
  lineBuffer_209 = _RAND_216[7:0];
  _RAND_217 = {1{`RANDOM}};
  lineBuffer_210 = _RAND_217[7:0];
  _RAND_218 = {1{`RANDOM}};
  lineBuffer_211 = _RAND_218[7:0];
  _RAND_219 = {1{`RANDOM}};
  lineBuffer_212 = _RAND_219[7:0];
  _RAND_220 = {1{`RANDOM}};
  lineBuffer_213 = _RAND_220[7:0];
  _RAND_221 = {1{`RANDOM}};
  lineBuffer_214 = _RAND_221[7:0];
  _RAND_222 = {1{`RANDOM}};
  lineBuffer_215 = _RAND_222[7:0];
  _RAND_223 = {1{`RANDOM}};
  lineBuffer_216 = _RAND_223[7:0];
  _RAND_224 = {1{`RANDOM}};
  lineBuffer_217 = _RAND_224[7:0];
  _RAND_225 = {1{`RANDOM}};
  lineBuffer_218 = _RAND_225[7:0];
  _RAND_226 = {1{`RANDOM}};
  lineBuffer_219 = _RAND_226[7:0];
  _RAND_227 = {1{`RANDOM}};
  lineBuffer_220 = _RAND_227[7:0];
  _RAND_228 = {1{`RANDOM}};
  lineBuffer_221 = _RAND_228[7:0];
  _RAND_229 = {1{`RANDOM}};
  lineBuffer_222 = _RAND_229[7:0];
  _RAND_230 = {1{`RANDOM}};
  lineBuffer_223 = _RAND_230[7:0];
  _RAND_231 = {1{`RANDOM}};
  lineBuffer_224 = _RAND_231[7:0];
  _RAND_232 = {1{`RANDOM}};
  lineBuffer_225 = _RAND_232[7:0];
  _RAND_233 = {1{`RANDOM}};
  lineBuffer_226 = _RAND_233[7:0];
  _RAND_234 = {1{`RANDOM}};
  lineBuffer_227 = _RAND_234[7:0];
  _RAND_235 = {1{`RANDOM}};
  lineBuffer_228 = _RAND_235[7:0];
  _RAND_236 = {1{`RANDOM}};
  lineBuffer_229 = _RAND_236[7:0];
  _RAND_237 = {1{`RANDOM}};
  lineBuffer_230 = _RAND_237[7:0];
  _RAND_238 = {1{`RANDOM}};
  lineBuffer_231 = _RAND_238[7:0];
  _RAND_239 = {1{`RANDOM}};
  lineBuffer_232 = _RAND_239[7:0];
  _RAND_240 = {1{`RANDOM}};
  lineBuffer_233 = _RAND_240[7:0];
  _RAND_241 = {1{`RANDOM}};
  lineBuffer_234 = _RAND_241[7:0];
  _RAND_242 = {1{`RANDOM}};
  lineBuffer_235 = _RAND_242[7:0];
  _RAND_243 = {1{`RANDOM}};
  lineBuffer_236 = _RAND_243[7:0];
  _RAND_244 = {1{`RANDOM}};
  lineBuffer_237 = _RAND_244[7:0];
  _RAND_245 = {1{`RANDOM}};
  lineBuffer_238 = _RAND_245[7:0];
  _RAND_246 = {1{`RANDOM}};
  lineBuffer_239 = _RAND_246[7:0];
  _RAND_247 = {1{`RANDOM}};
  lineBuffer_240 = _RAND_247[7:0];
  _RAND_248 = {1{`RANDOM}};
  lineBuffer_241 = _RAND_248[7:0];
  _RAND_249 = {1{`RANDOM}};
  lineBuffer_242 = _RAND_249[7:0];
  _RAND_250 = {1{`RANDOM}};
  lineBuffer_243 = _RAND_250[7:0];
  _RAND_251 = {1{`RANDOM}};
  lineBuffer_244 = _RAND_251[7:0];
  _RAND_252 = {1{`RANDOM}};
  lineBuffer_245 = _RAND_252[7:0];
  _RAND_253 = {1{`RANDOM}};
  lineBuffer_246 = _RAND_253[7:0];
  _RAND_254 = {1{`RANDOM}};
  lineBuffer_247 = _RAND_254[7:0];
  _RAND_255 = {1{`RANDOM}};
  lineBuffer_248 = _RAND_255[7:0];
  _RAND_256 = {1{`RANDOM}};
  lineBuffer_249 = _RAND_256[7:0];
  _RAND_257 = {1{`RANDOM}};
  lineBuffer_250 = _RAND_257[7:0];
  _RAND_258 = {1{`RANDOM}};
  lineBuffer_251 = _RAND_258[7:0];
  _RAND_259 = {1{`RANDOM}};
  lineBuffer_252 = _RAND_259[7:0];
  _RAND_260 = {1{`RANDOM}};
  lineBuffer_253 = _RAND_260[7:0];
  _RAND_261 = {1{`RANDOM}};
  lineBuffer_254 = _RAND_261[7:0];
  _RAND_262 = {1{`RANDOM}};
  lineBuffer_255 = _RAND_262[7:0];
  _RAND_263 = {1{`RANDOM}};
  lineBuffer_256 = _RAND_263[7:0];
  _RAND_264 = {1{`RANDOM}};
  lineBuffer_257 = _RAND_264[7:0];
  _RAND_265 = {1{`RANDOM}};
  lineBuffer_258 = _RAND_265[7:0];
  _RAND_266 = {1{`RANDOM}};
  lineBuffer_259 = _RAND_266[7:0];
  _RAND_267 = {1{`RANDOM}};
  lineBuffer_260 = _RAND_267[7:0];
  _RAND_268 = {1{`RANDOM}};
  lineBuffer_261 = _RAND_268[7:0];
  _RAND_269 = {1{`RANDOM}};
  lineBuffer_262 = _RAND_269[7:0];
  _RAND_270 = {1{`RANDOM}};
  lineBuffer_263 = _RAND_270[7:0];
  _RAND_271 = {1{`RANDOM}};
  lineBuffer_264 = _RAND_271[7:0];
  _RAND_272 = {1{`RANDOM}};
  lineBuffer_265 = _RAND_272[7:0];
  _RAND_273 = {1{`RANDOM}};
  lineBuffer_266 = _RAND_273[7:0];
  _RAND_274 = {1{`RANDOM}};
  lineBuffer_267 = _RAND_274[7:0];
  _RAND_275 = {1{`RANDOM}};
  lineBuffer_268 = _RAND_275[7:0];
  _RAND_276 = {1{`RANDOM}};
  lineBuffer_269 = _RAND_276[7:0];
  _RAND_277 = {1{`RANDOM}};
  lineBuffer_270 = _RAND_277[7:0];
  _RAND_278 = {1{`RANDOM}};
  lineBuffer_271 = _RAND_278[7:0];
  _RAND_279 = {1{`RANDOM}};
  lineBuffer_272 = _RAND_279[7:0];
  _RAND_280 = {1{`RANDOM}};
  lineBuffer_273 = _RAND_280[7:0];
  _RAND_281 = {1{`RANDOM}};
  lineBuffer_274 = _RAND_281[7:0];
  _RAND_282 = {1{`RANDOM}};
  lineBuffer_275 = _RAND_282[7:0];
  _RAND_283 = {1{`RANDOM}};
  lineBuffer_276 = _RAND_283[7:0];
  _RAND_284 = {1{`RANDOM}};
  lineBuffer_277 = _RAND_284[7:0];
  _RAND_285 = {1{`RANDOM}};
  lineBuffer_278 = _RAND_285[7:0];
  _RAND_286 = {1{`RANDOM}};
  lineBuffer_279 = _RAND_286[7:0];
  _RAND_287 = {1{`RANDOM}};
  lineBuffer_280 = _RAND_287[7:0];
  _RAND_288 = {1{`RANDOM}};
  lineBuffer_281 = _RAND_288[7:0];
  _RAND_289 = {1{`RANDOM}};
  lineBuffer_282 = _RAND_289[7:0];
  _RAND_290 = {1{`RANDOM}};
  lineBuffer_283 = _RAND_290[7:0];
  _RAND_291 = {1{`RANDOM}};
  lineBuffer_284 = _RAND_291[7:0];
  _RAND_292 = {1{`RANDOM}};
  lineBuffer_285 = _RAND_292[7:0];
  _RAND_293 = {1{`RANDOM}};
  lineBuffer_286 = _RAND_293[7:0];
  _RAND_294 = {1{`RANDOM}};
  lineBuffer_287 = _RAND_294[7:0];
  _RAND_295 = {1{`RANDOM}};
  lineBuffer_288 = _RAND_295[7:0];
  _RAND_296 = {1{`RANDOM}};
  lineBuffer_289 = _RAND_296[7:0];
  _RAND_297 = {1{`RANDOM}};
  lineBuffer_290 = _RAND_297[7:0];
  _RAND_298 = {1{`RANDOM}};
  lineBuffer_291 = _RAND_298[7:0];
  _RAND_299 = {1{`RANDOM}};
  lineBuffer_292 = _RAND_299[7:0];
  _RAND_300 = {1{`RANDOM}};
  lineBuffer_293 = _RAND_300[7:0];
  _RAND_301 = {1{`RANDOM}};
  lineBuffer_294 = _RAND_301[7:0];
  _RAND_302 = {1{`RANDOM}};
  lineBuffer_295 = _RAND_302[7:0];
  _RAND_303 = {1{`RANDOM}};
  lineBuffer_296 = _RAND_303[7:0];
  _RAND_304 = {1{`RANDOM}};
  lineBuffer_297 = _RAND_304[7:0];
  _RAND_305 = {1{`RANDOM}};
  lineBuffer_298 = _RAND_305[7:0];
  _RAND_306 = {1{`RANDOM}};
  lineBuffer_299 = _RAND_306[7:0];
  _RAND_307 = {1{`RANDOM}};
  lineBuffer_300 = _RAND_307[7:0];
  _RAND_308 = {1{`RANDOM}};
  lineBuffer_301 = _RAND_308[7:0];
  _RAND_309 = {1{`RANDOM}};
  lineBuffer_302 = _RAND_309[7:0];
  _RAND_310 = {1{`RANDOM}};
  lineBuffer_303 = _RAND_310[7:0];
  _RAND_311 = {1{`RANDOM}};
  lineBuffer_304 = _RAND_311[7:0];
  _RAND_312 = {1{`RANDOM}};
  lineBuffer_305 = _RAND_312[7:0];
  _RAND_313 = {1{`RANDOM}};
  lineBuffer_306 = _RAND_313[7:0];
  _RAND_314 = {1{`RANDOM}};
  lineBuffer_307 = _RAND_314[7:0];
  _RAND_315 = {1{`RANDOM}};
  lineBuffer_308 = _RAND_315[7:0];
  _RAND_316 = {1{`RANDOM}};
  lineBuffer_309 = _RAND_316[7:0];
  _RAND_317 = {1{`RANDOM}};
  lineBuffer_310 = _RAND_317[7:0];
  _RAND_318 = {1{`RANDOM}};
  lineBuffer_311 = _RAND_318[7:0];
  _RAND_319 = {1{`RANDOM}};
  lineBuffer_312 = _RAND_319[7:0];
  _RAND_320 = {1{`RANDOM}};
  lineBuffer_313 = _RAND_320[7:0];
  _RAND_321 = {1{`RANDOM}};
  lineBuffer_314 = _RAND_321[7:0];
  _RAND_322 = {1{`RANDOM}};
  lineBuffer_315 = _RAND_322[7:0];
  _RAND_323 = {1{`RANDOM}};
  lineBuffer_316 = _RAND_323[7:0];
  _RAND_324 = {1{`RANDOM}};
  lineBuffer_317 = _RAND_324[7:0];
  _RAND_325 = {1{`RANDOM}};
  lineBuffer_318 = _RAND_325[7:0];
  _RAND_326 = {1{`RANDOM}};
  lineBuffer_319 = _RAND_326[7:0];
  _RAND_327 = {1{`RANDOM}};
  lineBuffer_320 = _RAND_327[7:0];
  _RAND_328 = {1{`RANDOM}};
  lineBuffer_321 = _RAND_328[7:0];
  _RAND_329 = {1{`RANDOM}};
  lineBuffer_322 = _RAND_329[7:0];
  _RAND_330 = {1{`RANDOM}};
  lineBuffer_323 = _RAND_330[7:0];
  _RAND_331 = {1{`RANDOM}};
  lineBuffer_324 = _RAND_331[7:0];
  _RAND_332 = {1{`RANDOM}};
  lineBuffer_325 = _RAND_332[7:0];
  _RAND_333 = {1{`RANDOM}};
  lineBuffer_326 = _RAND_333[7:0];
  _RAND_334 = {1{`RANDOM}};
  lineBuffer_327 = _RAND_334[7:0];
  _RAND_335 = {1{`RANDOM}};
  lineBuffer_328 = _RAND_335[7:0];
  _RAND_336 = {1{`RANDOM}};
  lineBuffer_329 = _RAND_336[7:0];
  _RAND_337 = {1{`RANDOM}};
  lineBuffer_330 = _RAND_337[7:0];
  _RAND_338 = {1{`RANDOM}};
  lineBuffer_331 = _RAND_338[7:0];
  _RAND_339 = {1{`RANDOM}};
  lineBuffer_332 = _RAND_339[7:0];
  _RAND_340 = {1{`RANDOM}};
  lineBuffer_333 = _RAND_340[7:0];
  _RAND_341 = {1{`RANDOM}};
  lineBuffer_334 = _RAND_341[7:0];
  _RAND_342 = {1{`RANDOM}};
  lineBuffer_335 = _RAND_342[7:0];
  _RAND_343 = {1{`RANDOM}};
  lineBuffer_336 = _RAND_343[7:0];
  _RAND_344 = {1{`RANDOM}};
  lineBuffer_337 = _RAND_344[7:0];
  _RAND_345 = {1{`RANDOM}};
  lineBuffer_338 = _RAND_345[7:0];
  _RAND_346 = {1{`RANDOM}};
  lineBuffer_339 = _RAND_346[7:0];
  _RAND_347 = {1{`RANDOM}};
  lineBuffer_340 = _RAND_347[7:0];
  _RAND_348 = {1{`RANDOM}};
  lineBuffer_341 = _RAND_348[7:0];
  _RAND_349 = {1{`RANDOM}};
  lineBuffer_342 = _RAND_349[7:0];
  _RAND_350 = {1{`RANDOM}};
  lineBuffer_343 = _RAND_350[7:0];
  _RAND_351 = {1{`RANDOM}};
  lineBuffer_344 = _RAND_351[7:0];
  _RAND_352 = {1{`RANDOM}};
  lineBuffer_345 = _RAND_352[7:0];
  _RAND_353 = {1{`RANDOM}};
  lineBuffer_346 = _RAND_353[7:0];
  _RAND_354 = {1{`RANDOM}};
  lineBuffer_347 = _RAND_354[7:0];
  _RAND_355 = {1{`RANDOM}};
  lineBuffer_348 = _RAND_355[7:0];
  _RAND_356 = {1{`RANDOM}};
  lineBuffer_349 = _RAND_356[7:0];
  _RAND_357 = {1{`RANDOM}};
  lineBuffer_350 = _RAND_357[7:0];
  _RAND_358 = {1{`RANDOM}};
  lineBuffer_351 = _RAND_358[7:0];
  _RAND_359 = {1{`RANDOM}};
  lineBuffer_352 = _RAND_359[7:0];
  _RAND_360 = {1{`RANDOM}};
  lineBuffer_353 = _RAND_360[7:0];
  _RAND_361 = {1{`RANDOM}};
  lineBuffer_354 = _RAND_361[7:0];
  _RAND_362 = {1{`RANDOM}};
  lineBuffer_355 = _RAND_362[7:0];
  _RAND_363 = {1{`RANDOM}};
  lineBuffer_356 = _RAND_363[7:0];
  _RAND_364 = {1{`RANDOM}};
  lineBuffer_357 = _RAND_364[7:0];
  _RAND_365 = {1{`RANDOM}};
  lineBuffer_358 = _RAND_365[7:0];
  _RAND_366 = {1{`RANDOM}};
  lineBuffer_359 = _RAND_366[7:0];
  _RAND_367 = {1{`RANDOM}};
  lineBuffer_360 = _RAND_367[7:0];
  _RAND_368 = {1{`RANDOM}};
  lineBuffer_361 = _RAND_368[7:0];
  _RAND_369 = {1{`RANDOM}};
  lineBuffer_362 = _RAND_369[7:0];
  _RAND_370 = {1{`RANDOM}};
  lineBuffer_363 = _RAND_370[7:0];
  _RAND_371 = {1{`RANDOM}};
  lineBuffer_364 = _RAND_371[7:0];
  _RAND_372 = {1{`RANDOM}};
  lineBuffer_365 = _RAND_372[7:0];
  _RAND_373 = {1{`RANDOM}};
  lineBuffer_366 = _RAND_373[7:0];
  _RAND_374 = {1{`RANDOM}};
  lineBuffer_367 = _RAND_374[7:0];
  _RAND_375 = {1{`RANDOM}};
  lineBuffer_368 = _RAND_375[7:0];
  _RAND_376 = {1{`RANDOM}};
  lineBuffer_369 = _RAND_376[7:0];
  _RAND_377 = {1{`RANDOM}};
  lineBuffer_370 = _RAND_377[7:0];
  _RAND_378 = {1{`RANDOM}};
  lineBuffer_371 = _RAND_378[7:0];
  _RAND_379 = {1{`RANDOM}};
  lineBuffer_372 = _RAND_379[7:0];
  _RAND_380 = {1{`RANDOM}};
  lineBuffer_373 = _RAND_380[7:0];
  _RAND_381 = {1{`RANDOM}};
  lineBuffer_374 = _RAND_381[7:0];
  _RAND_382 = {1{`RANDOM}};
  lineBuffer_375 = _RAND_382[7:0];
  _RAND_383 = {1{`RANDOM}};
  lineBuffer_376 = _RAND_383[7:0];
  _RAND_384 = {1{`RANDOM}};
  lineBuffer_377 = _RAND_384[7:0];
  _RAND_385 = {1{`RANDOM}};
  lineBuffer_378 = _RAND_385[7:0];
  _RAND_386 = {1{`RANDOM}};
  lineBuffer_379 = _RAND_386[7:0];
  _RAND_387 = {1{`RANDOM}};
  lineBuffer_380 = _RAND_387[7:0];
  _RAND_388 = {1{`RANDOM}};
  lineBuffer_381 = _RAND_388[7:0];
  _RAND_389 = {1{`RANDOM}};
  lineBuffer_382 = _RAND_389[7:0];
  _RAND_390 = {1{`RANDOM}};
  lineBuffer_383 = _RAND_390[7:0];
  _RAND_391 = {1{`RANDOM}};
  lineBuffer_384 = _RAND_391[7:0];
  _RAND_392 = {1{`RANDOM}};
  lineBuffer_385 = _RAND_392[7:0];
  _RAND_393 = {1{`RANDOM}};
  lineBuffer_386 = _RAND_393[7:0];
  _RAND_394 = {1{`RANDOM}};
  lineBuffer_387 = _RAND_394[7:0];
  _RAND_395 = {1{`RANDOM}};
  lineBuffer_388 = _RAND_395[7:0];
  _RAND_396 = {1{`RANDOM}};
  lineBuffer_389 = _RAND_396[7:0];
  _RAND_397 = {1{`RANDOM}};
  lineBuffer_390 = _RAND_397[7:0];
  _RAND_398 = {1{`RANDOM}};
  lineBuffer_391 = _RAND_398[7:0];
  _RAND_399 = {1{`RANDOM}};
  lineBuffer_392 = _RAND_399[7:0];
  _RAND_400 = {1{`RANDOM}};
  lineBuffer_393 = _RAND_400[7:0];
  _RAND_401 = {1{`RANDOM}};
  lineBuffer_394 = _RAND_401[7:0];
  _RAND_402 = {1{`RANDOM}};
  lineBuffer_395 = _RAND_402[7:0];
  _RAND_403 = {1{`RANDOM}};
  lineBuffer_396 = _RAND_403[7:0];
  _RAND_404 = {1{`RANDOM}};
  lineBuffer_397 = _RAND_404[7:0];
  _RAND_405 = {1{`RANDOM}};
  lineBuffer_398 = _RAND_405[7:0];
  _RAND_406 = {1{`RANDOM}};
  lineBuffer_399 = _RAND_406[7:0];
  _RAND_407 = {1{`RANDOM}};
  lineBuffer_400 = _RAND_407[7:0];
  _RAND_408 = {1{`RANDOM}};
  lineBuffer_401 = _RAND_408[7:0];
  _RAND_409 = {1{`RANDOM}};
  lineBuffer_402 = _RAND_409[7:0];
  _RAND_410 = {1{`RANDOM}};
  lineBuffer_403 = _RAND_410[7:0];
  _RAND_411 = {1{`RANDOM}};
  lineBuffer_404 = _RAND_411[7:0];
  _RAND_412 = {1{`RANDOM}};
  lineBuffer_405 = _RAND_412[7:0];
  _RAND_413 = {1{`RANDOM}};
  lineBuffer_406 = _RAND_413[7:0];
  _RAND_414 = {1{`RANDOM}};
  lineBuffer_407 = _RAND_414[7:0];
  _RAND_415 = {1{`RANDOM}};
  lineBuffer_408 = _RAND_415[7:0];
  _RAND_416 = {1{`RANDOM}};
  lineBuffer_409 = _RAND_416[7:0];
  _RAND_417 = {1{`RANDOM}};
  lineBuffer_410 = _RAND_417[7:0];
  _RAND_418 = {1{`RANDOM}};
  lineBuffer_411 = _RAND_418[7:0];
  _RAND_419 = {1{`RANDOM}};
  lineBuffer_412 = _RAND_419[7:0];
  _RAND_420 = {1{`RANDOM}};
  lineBuffer_413 = _RAND_420[7:0];
  _RAND_421 = {1{`RANDOM}};
  lineBuffer_414 = _RAND_421[7:0];
  _RAND_422 = {1{`RANDOM}};
  lineBuffer_415 = _RAND_422[7:0];
  _RAND_423 = {1{`RANDOM}};
  lineBuffer_416 = _RAND_423[7:0];
  _RAND_424 = {1{`RANDOM}};
  lineBuffer_417 = _RAND_424[7:0];
  _RAND_425 = {1{`RANDOM}};
  lineBuffer_418 = _RAND_425[7:0];
  _RAND_426 = {1{`RANDOM}};
  lineBuffer_419 = _RAND_426[7:0];
  _RAND_427 = {1{`RANDOM}};
  lineBuffer_420 = _RAND_427[7:0];
  _RAND_428 = {1{`RANDOM}};
  lineBuffer_421 = _RAND_428[7:0];
  _RAND_429 = {1{`RANDOM}};
  lineBuffer_422 = _RAND_429[7:0];
  _RAND_430 = {1{`RANDOM}};
  lineBuffer_423 = _RAND_430[7:0];
  _RAND_431 = {1{`RANDOM}};
  lineBuffer_424 = _RAND_431[7:0];
  _RAND_432 = {1{`RANDOM}};
  lineBuffer_425 = _RAND_432[7:0];
  _RAND_433 = {1{`RANDOM}};
  lineBuffer_426 = _RAND_433[7:0];
  _RAND_434 = {1{`RANDOM}};
  lineBuffer_427 = _RAND_434[7:0];
  _RAND_435 = {1{`RANDOM}};
  lineBuffer_428 = _RAND_435[7:0];
  _RAND_436 = {1{`RANDOM}};
  lineBuffer_429 = _RAND_436[7:0];
  _RAND_437 = {1{`RANDOM}};
  lineBuffer_430 = _RAND_437[7:0];
  _RAND_438 = {1{`RANDOM}};
  lineBuffer_431 = _RAND_438[7:0];
  _RAND_439 = {1{`RANDOM}};
  lineBuffer_432 = _RAND_439[7:0];
  _RAND_440 = {1{`RANDOM}};
  lineBuffer_433 = _RAND_440[7:0];
  _RAND_441 = {1{`RANDOM}};
  lineBuffer_434 = _RAND_441[7:0];
  _RAND_442 = {1{`RANDOM}};
  lineBuffer_435 = _RAND_442[7:0];
  _RAND_443 = {1{`RANDOM}};
  lineBuffer_436 = _RAND_443[7:0];
  _RAND_444 = {1{`RANDOM}};
  lineBuffer_437 = _RAND_444[7:0];
  _RAND_445 = {1{`RANDOM}};
  lineBuffer_438 = _RAND_445[7:0];
  _RAND_446 = {1{`RANDOM}};
  lineBuffer_439 = _RAND_446[7:0];
  _RAND_447 = {1{`RANDOM}};
  lineBuffer_440 = _RAND_447[7:0];
  _RAND_448 = {1{`RANDOM}};
  lineBuffer_441 = _RAND_448[7:0];
  _RAND_449 = {1{`RANDOM}};
  lineBuffer_442 = _RAND_449[7:0];
  _RAND_450 = {1{`RANDOM}};
  lineBuffer_443 = _RAND_450[7:0];
  _RAND_451 = {1{`RANDOM}};
  lineBuffer_444 = _RAND_451[7:0];
  _RAND_452 = {1{`RANDOM}};
  lineBuffer_445 = _RAND_452[7:0];
  _RAND_453 = {1{`RANDOM}};
  lineBuffer_446 = _RAND_453[7:0];
  _RAND_454 = {1{`RANDOM}};
  lineBuffer_447 = _RAND_454[7:0];
  _RAND_455 = {1{`RANDOM}};
  lineBuffer_448 = _RAND_455[7:0];
  _RAND_456 = {1{`RANDOM}};
  lineBuffer_449 = _RAND_456[7:0];
  _RAND_457 = {1{`RANDOM}};
  lineBuffer_450 = _RAND_457[7:0];
  _RAND_458 = {1{`RANDOM}};
  lineBuffer_451 = _RAND_458[7:0];
  _RAND_459 = {1{`RANDOM}};
  lineBuffer_452 = _RAND_459[7:0];
  _RAND_460 = {1{`RANDOM}};
  lineBuffer_453 = _RAND_460[7:0];
  _RAND_461 = {1{`RANDOM}};
  lineBuffer_454 = _RAND_461[7:0];
  _RAND_462 = {1{`RANDOM}};
  lineBuffer_455 = _RAND_462[7:0];
  _RAND_463 = {1{`RANDOM}};
  lineBuffer_456 = _RAND_463[7:0];
  _RAND_464 = {1{`RANDOM}};
  lineBuffer_457 = _RAND_464[7:0];
  _RAND_465 = {1{`RANDOM}};
  lineBuffer_458 = _RAND_465[7:0];
  _RAND_466 = {1{`RANDOM}};
  lineBuffer_459 = _RAND_466[7:0];
  _RAND_467 = {1{`RANDOM}};
  lineBuffer_460 = _RAND_467[7:0];
  _RAND_468 = {1{`RANDOM}};
  lineBuffer_461 = _RAND_468[7:0];
  _RAND_469 = {1{`RANDOM}};
  lineBuffer_462 = _RAND_469[7:0];
  _RAND_470 = {1{`RANDOM}};
  lineBuffer_463 = _RAND_470[7:0];
  _RAND_471 = {1{`RANDOM}};
  lineBuffer_464 = _RAND_471[7:0];
  _RAND_472 = {1{`RANDOM}};
  lineBuffer_465 = _RAND_472[7:0];
  _RAND_473 = {1{`RANDOM}};
  lineBuffer_466 = _RAND_473[7:0];
  _RAND_474 = {1{`RANDOM}};
  lineBuffer_467 = _RAND_474[7:0];
  _RAND_475 = {1{`RANDOM}};
  lineBuffer_468 = _RAND_475[7:0];
  _RAND_476 = {1{`RANDOM}};
  lineBuffer_469 = _RAND_476[7:0];
  _RAND_477 = {1{`RANDOM}};
  lineBuffer_470 = _RAND_477[7:0];
  _RAND_478 = {1{`RANDOM}};
  lineBuffer_471 = _RAND_478[7:0];
  _RAND_479 = {1{`RANDOM}};
  lineBuffer_472 = _RAND_479[7:0];
  _RAND_480 = {1{`RANDOM}};
  lineBuffer_473 = _RAND_480[7:0];
  _RAND_481 = {1{`RANDOM}};
  lineBuffer_474 = _RAND_481[7:0];
  _RAND_482 = {1{`RANDOM}};
  lineBuffer_475 = _RAND_482[7:0];
  _RAND_483 = {1{`RANDOM}};
  lineBuffer_476 = _RAND_483[7:0];
  _RAND_484 = {1{`RANDOM}};
  lineBuffer_477 = _RAND_484[7:0];
  _RAND_485 = {1{`RANDOM}};
  lineBuffer_478 = _RAND_485[7:0];
  _RAND_486 = {1{`RANDOM}};
  lineBuffer_479 = _RAND_486[7:0];
  _RAND_487 = {1{`RANDOM}};
  lineBuffer_480 = _RAND_487[7:0];
  _RAND_488 = {1{`RANDOM}};
  lineBuffer_481 = _RAND_488[7:0];
  _RAND_489 = {1{`RANDOM}};
  lineBuffer_482 = _RAND_489[7:0];
  _RAND_490 = {1{`RANDOM}};
  lineBuffer_483 = _RAND_490[7:0];
  _RAND_491 = {1{`RANDOM}};
  lineBuffer_484 = _RAND_491[7:0];
  _RAND_492 = {1{`RANDOM}};
  lineBuffer_485 = _RAND_492[7:0];
  _RAND_493 = {1{`RANDOM}};
  lineBuffer_486 = _RAND_493[7:0];
  _RAND_494 = {1{`RANDOM}};
  lineBuffer_487 = _RAND_494[7:0];
  _RAND_495 = {1{`RANDOM}};
  lineBuffer_488 = _RAND_495[7:0];
  _RAND_496 = {1{`RANDOM}};
  lineBuffer_489 = _RAND_496[7:0];
  _RAND_497 = {1{`RANDOM}};
  lineBuffer_490 = _RAND_497[7:0];
  _RAND_498 = {1{`RANDOM}};
  lineBuffer_491 = _RAND_498[7:0];
  _RAND_499 = {1{`RANDOM}};
  lineBuffer_492 = _RAND_499[7:0];
  _RAND_500 = {1{`RANDOM}};
  lineBuffer_493 = _RAND_500[7:0];
  _RAND_501 = {1{`RANDOM}};
  lineBuffer_494 = _RAND_501[7:0];
  _RAND_502 = {1{`RANDOM}};
  lineBuffer_495 = _RAND_502[7:0];
  _RAND_503 = {1{`RANDOM}};
  lineBuffer_496 = _RAND_503[7:0];
  _RAND_504 = {1{`RANDOM}};
  lineBuffer_497 = _RAND_504[7:0];
  _RAND_505 = {1{`RANDOM}};
  lineBuffer_498 = _RAND_505[7:0];
  _RAND_506 = {1{`RANDOM}};
  lineBuffer_499 = _RAND_506[7:0];
  _RAND_507 = {1{`RANDOM}};
  lineBuffer_500 = _RAND_507[7:0];
  _RAND_508 = {1{`RANDOM}};
  lineBuffer_501 = _RAND_508[7:0];
  _RAND_509 = {1{`RANDOM}};
  lineBuffer_502 = _RAND_509[7:0];
  _RAND_510 = {1{`RANDOM}};
  lineBuffer_503 = _RAND_510[7:0];
  _RAND_511 = {1{`RANDOM}};
  lineBuffer_504 = _RAND_511[7:0];
  _RAND_512 = {1{`RANDOM}};
  lineBuffer_505 = _RAND_512[7:0];
  _RAND_513 = {1{`RANDOM}};
  lineBuffer_506 = _RAND_513[7:0];
  _RAND_514 = {1{`RANDOM}};
  lineBuffer_507 = _RAND_514[7:0];
  _RAND_515 = {1{`RANDOM}};
  lineBuffer_508 = _RAND_515[7:0];
  _RAND_516 = {1{`RANDOM}};
  lineBuffer_509 = _RAND_516[7:0];
  _RAND_517 = {1{`RANDOM}};
  lineBuffer_510 = _RAND_517[7:0];
  _RAND_518 = {1{`RANDOM}};
  lineBuffer_511 = _RAND_518[7:0];
  _RAND_519 = {1{`RANDOM}};
  lineBuffer_512 = _RAND_519[7:0];
  _RAND_520 = {1{`RANDOM}};
  lineBuffer_513 = _RAND_520[7:0];
  _RAND_521 = {1{`RANDOM}};
  lineBuffer_514 = _RAND_521[7:0];
  _RAND_522 = {1{`RANDOM}};
  lineBuffer_515 = _RAND_522[7:0];
  _RAND_523 = {1{`RANDOM}};
  lineBuffer_516 = _RAND_523[7:0];
  _RAND_524 = {1{`RANDOM}};
  lineBuffer_517 = _RAND_524[7:0];
  _RAND_525 = {1{`RANDOM}};
  lineBuffer_518 = _RAND_525[7:0];
  _RAND_526 = {1{`RANDOM}};
  lineBuffer_519 = _RAND_526[7:0];
  _RAND_527 = {1{`RANDOM}};
  lineBuffer_520 = _RAND_527[7:0];
  _RAND_528 = {1{`RANDOM}};
  lineBuffer_521 = _RAND_528[7:0];
  _RAND_529 = {1{`RANDOM}};
  lineBuffer_522 = _RAND_529[7:0];
  _RAND_530 = {1{`RANDOM}};
  lineBuffer_523 = _RAND_530[7:0];
  _RAND_531 = {1{`RANDOM}};
  lineBuffer_524 = _RAND_531[7:0];
  _RAND_532 = {1{`RANDOM}};
  lineBuffer_525 = _RAND_532[7:0];
  _RAND_533 = {1{`RANDOM}};
  lineBuffer_526 = _RAND_533[7:0];
  _RAND_534 = {1{`RANDOM}};
  lineBuffer_527 = _RAND_534[7:0];
  _RAND_535 = {1{`RANDOM}};
  lineBuffer_528 = _RAND_535[7:0];
  _RAND_536 = {1{`RANDOM}};
  lineBuffer_529 = _RAND_536[7:0];
  _RAND_537 = {1{`RANDOM}};
  lineBuffer_530 = _RAND_537[7:0];
  _RAND_538 = {1{`RANDOM}};
  lineBuffer_531 = _RAND_538[7:0];
  _RAND_539 = {1{`RANDOM}};
  lineBuffer_532 = _RAND_539[7:0];
  _RAND_540 = {1{`RANDOM}};
  lineBuffer_533 = _RAND_540[7:0];
  _RAND_541 = {1{`RANDOM}};
  lineBuffer_534 = _RAND_541[7:0];
  _RAND_542 = {1{`RANDOM}};
  lineBuffer_535 = _RAND_542[7:0];
  _RAND_543 = {1{`RANDOM}};
  lineBuffer_536 = _RAND_543[7:0];
  _RAND_544 = {1{`RANDOM}};
  lineBuffer_537 = _RAND_544[7:0];
  _RAND_545 = {1{`RANDOM}};
  lineBuffer_538 = _RAND_545[7:0];
  _RAND_546 = {1{`RANDOM}};
  lineBuffer_539 = _RAND_546[7:0];
  _RAND_547 = {1{`RANDOM}};
  lineBuffer_540 = _RAND_547[7:0];
  _RAND_548 = {1{`RANDOM}};
  lineBuffer_541 = _RAND_548[7:0];
  _RAND_549 = {1{`RANDOM}};
  lineBuffer_542 = _RAND_549[7:0];
  _RAND_550 = {1{`RANDOM}};
  lineBuffer_543 = _RAND_550[7:0];
  _RAND_551 = {1{`RANDOM}};
  lineBuffer_544 = _RAND_551[7:0];
  _RAND_552 = {1{`RANDOM}};
  lineBuffer_545 = _RAND_552[7:0];
  _RAND_553 = {1{`RANDOM}};
  lineBuffer_546 = _RAND_553[7:0];
  _RAND_554 = {1{`RANDOM}};
  lineBuffer_547 = _RAND_554[7:0];
  _RAND_555 = {1{`RANDOM}};
  lineBuffer_548 = _RAND_555[7:0];
  _RAND_556 = {1{`RANDOM}};
  lineBuffer_549 = _RAND_556[7:0];
  _RAND_557 = {1{`RANDOM}};
  lineBuffer_550 = _RAND_557[7:0];
  _RAND_558 = {1{`RANDOM}};
  lineBuffer_551 = _RAND_558[7:0];
  _RAND_559 = {1{`RANDOM}};
  lineBuffer_552 = _RAND_559[7:0];
  _RAND_560 = {1{`RANDOM}};
  lineBuffer_553 = _RAND_560[7:0];
  _RAND_561 = {1{`RANDOM}};
  lineBuffer_554 = _RAND_561[7:0];
  _RAND_562 = {1{`RANDOM}};
  lineBuffer_555 = _RAND_562[7:0];
  _RAND_563 = {1{`RANDOM}};
  lineBuffer_556 = _RAND_563[7:0];
  _RAND_564 = {1{`RANDOM}};
  lineBuffer_557 = _RAND_564[7:0];
  _RAND_565 = {1{`RANDOM}};
  lineBuffer_558 = _RAND_565[7:0];
  _RAND_566 = {1{`RANDOM}};
  lineBuffer_559 = _RAND_566[7:0];
  _RAND_567 = {1{`RANDOM}};
  lineBuffer_560 = _RAND_567[7:0];
  _RAND_568 = {1{`RANDOM}};
  lineBuffer_561 = _RAND_568[7:0];
  _RAND_569 = {1{`RANDOM}};
  lineBuffer_562 = _RAND_569[7:0];
  _RAND_570 = {1{`RANDOM}};
  lineBuffer_563 = _RAND_570[7:0];
  _RAND_571 = {1{`RANDOM}};
  lineBuffer_564 = _RAND_571[7:0];
  _RAND_572 = {1{`RANDOM}};
  lineBuffer_565 = _RAND_572[7:0];
  _RAND_573 = {1{`RANDOM}};
  lineBuffer_566 = _RAND_573[7:0];
  _RAND_574 = {1{`RANDOM}};
  lineBuffer_567 = _RAND_574[7:0];
  _RAND_575 = {1{`RANDOM}};
  lineBuffer_568 = _RAND_575[7:0];
  _RAND_576 = {1{`RANDOM}};
  lineBuffer_569 = _RAND_576[7:0];
  _RAND_577 = {1{`RANDOM}};
  lineBuffer_570 = _RAND_577[7:0];
  _RAND_578 = {1{`RANDOM}};
  lineBuffer_571 = _RAND_578[7:0];
  _RAND_579 = {1{`RANDOM}};
  lineBuffer_572 = _RAND_579[7:0];
  _RAND_580 = {1{`RANDOM}};
  lineBuffer_573 = _RAND_580[7:0];
  _RAND_581 = {1{`RANDOM}};
  lineBuffer_574 = _RAND_581[7:0];
  _RAND_582 = {1{`RANDOM}};
  lineBuffer_575 = _RAND_582[7:0];
  _RAND_583 = {1{`RANDOM}};
  lineBuffer_576 = _RAND_583[7:0];
  _RAND_584 = {1{`RANDOM}};
  lineBuffer_577 = _RAND_584[7:0];
  _RAND_585 = {1{`RANDOM}};
  lineBuffer_578 = _RAND_585[7:0];
  _RAND_586 = {1{`RANDOM}};
  lineBuffer_579 = _RAND_586[7:0];
  _RAND_587 = {1{`RANDOM}};
  lineBuffer_580 = _RAND_587[7:0];
  _RAND_588 = {1{`RANDOM}};
  lineBuffer_581 = _RAND_588[7:0];
  _RAND_589 = {1{`RANDOM}};
  lineBuffer_582 = _RAND_589[7:0];
  _RAND_590 = {1{`RANDOM}};
  lineBuffer_583 = _RAND_590[7:0];
  _RAND_591 = {1{`RANDOM}};
  lineBuffer_584 = _RAND_591[7:0];
  _RAND_592 = {1{`RANDOM}};
  lineBuffer_585 = _RAND_592[7:0];
  _RAND_593 = {1{`RANDOM}};
  lineBuffer_586 = _RAND_593[7:0];
  _RAND_594 = {1{`RANDOM}};
  lineBuffer_587 = _RAND_594[7:0];
  _RAND_595 = {1{`RANDOM}};
  lineBuffer_588 = _RAND_595[7:0];
  _RAND_596 = {1{`RANDOM}};
  lineBuffer_589 = _RAND_596[7:0];
  _RAND_597 = {1{`RANDOM}};
  lineBuffer_590 = _RAND_597[7:0];
  _RAND_598 = {1{`RANDOM}};
  lineBuffer_591 = _RAND_598[7:0];
  _RAND_599 = {1{`RANDOM}};
  lineBuffer_592 = _RAND_599[7:0];
  _RAND_600 = {1{`RANDOM}};
  lineBuffer_593 = _RAND_600[7:0];
  _RAND_601 = {1{`RANDOM}};
  lineBuffer_594 = _RAND_601[7:0];
  _RAND_602 = {1{`RANDOM}};
  lineBuffer_595 = _RAND_602[7:0];
  _RAND_603 = {1{`RANDOM}};
  lineBuffer_596 = _RAND_603[7:0];
  _RAND_604 = {1{`RANDOM}};
  lineBuffer_597 = _RAND_604[7:0];
  _RAND_605 = {1{`RANDOM}};
  lineBuffer_598 = _RAND_605[7:0];
  _RAND_606 = {1{`RANDOM}};
  lineBuffer_599 = _RAND_606[7:0];
  _RAND_607 = {1{`RANDOM}};
  lineBuffer_600 = _RAND_607[7:0];
  _RAND_608 = {1{`RANDOM}};
  lineBuffer_601 = _RAND_608[7:0];
  _RAND_609 = {1{`RANDOM}};
  lineBuffer_602 = _RAND_609[7:0];
  _RAND_610 = {1{`RANDOM}};
  lineBuffer_603 = _RAND_610[7:0];
  _RAND_611 = {1{`RANDOM}};
  lineBuffer_604 = _RAND_611[7:0];
  _RAND_612 = {1{`RANDOM}};
  lineBuffer_605 = _RAND_612[7:0];
  _RAND_613 = {1{`RANDOM}};
  lineBuffer_606 = _RAND_613[7:0];
  _RAND_614 = {1{`RANDOM}};
  lineBuffer_607 = _RAND_614[7:0];
  _RAND_615 = {1{`RANDOM}};
  lineBuffer_608 = _RAND_615[7:0];
  _RAND_616 = {1{`RANDOM}};
  lineBuffer_609 = _RAND_616[7:0];
  _RAND_617 = {1{`RANDOM}};
  lineBuffer_610 = _RAND_617[7:0];
  _RAND_618 = {1{`RANDOM}};
  lineBuffer_611 = _RAND_618[7:0];
  _RAND_619 = {1{`RANDOM}};
  lineBuffer_612 = _RAND_619[7:0];
  _RAND_620 = {1{`RANDOM}};
  lineBuffer_613 = _RAND_620[7:0];
  _RAND_621 = {1{`RANDOM}};
  lineBuffer_614 = _RAND_621[7:0];
  _RAND_622 = {1{`RANDOM}};
  lineBuffer_615 = _RAND_622[7:0];
  _RAND_623 = {1{`RANDOM}};
  lineBuffer_616 = _RAND_623[7:0];
  _RAND_624 = {1{`RANDOM}};
  lineBuffer_617 = _RAND_624[7:0];
  _RAND_625 = {1{`RANDOM}};
  lineBuffer_618 = _RAND_625[7:0];
  _RAND_626 = {1{`RANDOM}};
  lineBuffer_619 = _RAND_626[7:0];
  _RAND_627 = {1{`RANDOM}};
  lineBuffer_620 = _RAND_627[7:0];
  _RAND_628 = {1{`RANDOM}};
  lineBuffer_621 = _RAND_628[7:0];
  _RAND_629 = {1{`RANDOM}};
  lineBuffer_622 = _RAND_629[7:0];
  _RAND_630 = {1{`RANDOM}};
  lineBuffer_623 = _RAND_630[7:0];
  _RAND_631 = {1{`RANDOM}};
  lineBuffer_624 = _RAND_631[7:0];
  _RAND_632 = {1{`RANDOM}};
  lineBuffer_625 = _RAND_632[7:0];
  _RAND_633 = {1{`RANDOM}};
  lineBuffer_626 = _RAND_633[7:0];
  _RAND_634 = {1{`RANDOM}};
  lineBuffer_627 = _RAND_634[7:0];
  _RAND_635 = {1{`RANDOM}};
  lineBuffer_628 = _RAND_635[7:0];
  _RAND_636 = {1{`RANDOM}};
  lineBuffer_629 = _RAND_636[7:0];
  _RAND_637 = {1{`RANDOM}};
  lineBuffer_630 = _RAND_637[7:0];
  _RAND_638 = {1{`RANDOM}};
  lineBuffer_631 = _RAND_638[7:0];
  _RAND_639 = {1{`RANDOM}};
  lineBuffer_632 = _RAND_639[7:0];
  _RAND_640 = {1{`RANDOM}};
  lineBuffer_633 = _RAND_640[7:0];
  _RAND_641 = {1{`RANDOM}};
  lineBuffer_634 = _RAND_641[7:0];
  _RAND_642 = {1{`RANDOM}};
  lineBuffer_635 = _RAND_642[7:0];
  _RAND_643 = {1{`RANDOM}};
  lineBuffer_636 = _RAND_643[7:0];
  _RAND_644 = {1{`RANDOM}};
  lineBuffer_637 = _RAND_644[7:0];
  _RAND_645 = {1{`RANDOM}};
  lineBuffer_638 = _RAND_645[7:0];
  _RAND_646 = {1{`RANDOM}};
  lineBuffer_639 = _RAND_646[7:0];
  _RAND_647 = {1{`RANDOM}};
  lineBuffer_640 = _RAND_647[7:0];
  _RAND_648 = {1{`RANDOM}};
  lineBuffer_641 = _RAND_648[7:0];
  _RAND_649 = {1{`RANDOM}};
  lineBuffer_642 = _RAND_649[7:0];
  _RAND_650 = {1{`RANDOM}};
  lineBuffer_643 = _RAND_650[7:0];
  _RAND_651 = {1{`RANDOM}};
  lineBuffer_644 = _RAND_651[7:0];
  _RAND_652 = {1{`RANDOM}};
  lineBuffer_645 = _RAND_652[7:0];
  _RAND_653 = {1{`RANDOM}};
  lineBuffer_646 = _RAND_653[7:0];
  _RAND_654 = {1{`RANDOM}};
  lineBuffer_647 = _RAND_654[7:0];
  _RAND_655 = {1{`RANDOM}};
  lineBuffer_648 = _RAND_655[7:0];
  _RAND_656 = {1{`RANDOM}};
  lineBuffer_649 = _RAND_656[7:0];
  _RAND_657 = {1{`RANDOM}};
  lineBuffer_650 = _RAND_657[7:0];
  _RAND_658 = {1{`RANDOM}};
  lineBuffer_651 = _RAND_658[7:0];
  _RAND_659 = {1{`RANDOM}};
  lineBuffer_652 = _RAND_659[7:0];
  _RAND_660 = {1{`RANDOM}};
  lineBuffer_653 = _RAND_660[7:0];
  _RAND_661 = {1{`RANDOM}};
  lineBuffer_654 = _RAND_661[7:0];
  _RAND_662 = {1{`RANDOM}};
  lineBuffer_655 = _RAND_662[7:0];
  _RAND_663 = {1{`RANDOM}};
  lineBuffer_656 = _RAND_663[7:0];
  _RAND_664 = {1{`RANDOM}};
  lineBuffer_657 = _RAND_664[7:0];
  _RAND_665 = {1{`RANDOM}};
  lineBuffer_658 = _RAND_665[7:0];
  _RAND_666 = {1{`RANDOM}};
  lineBuffer_659 = _RAND_666[7:0];
  _RAND_667 = {1{`RANDOM}};
  lineBuffer_660 = _RAND_667[7:0];
  _RAND_668 = {1{`RANDOM}};
  lineBuffer_661 = _RAND_668[7:0];
  _RAND_669 = {1{`RANDOM}};
  lineBuffer_662 = _RAND_669[7:0];
  _RAND_670 = {1{`RANDOM}};
  lineBuffer_663 = _RAND_670[7:0];
  _RAND_671 = {1{`RANDOM}};
  lineBuffer_664 = _RAND_671[7:0];
  _RAND_672 = {1{`RANDOM}};
  lineBuffer_665 = _RAND_672[7:0];
  _RAND_673 = {1{`RANDOM}};
  lineBuffer_666 = _RAND_673[7:0];
  _RAND_674 = {1{`RANDOM}};
  lineBuffer_667 = _RAND_674[7:0];
  _RAND_675 = {1{`RANDOM}};
  lineBuffer_668 = _RAND_675[7:0];
  _RAND_676 = {1{`RANDOM}};
  lineBuffer_669 = _RAND_676[7:0];
  _RAND_677 = {1{`RANDOM}};
  lineBuffer_670 = _RAND_677[7:0];
  _RAND_678 = {1{`RANDOM}};
  lineBuffer_671 = _RAND_678[7:0];
  _RAND_679 = {1{`RANDOM}};
  lineBuffer_672 = _RAND_679[7:0];
  _RAND_680 = {1{`RANDOM}};
  lineBuffer_673 = _RAND_680[7:0];
  _RAND_681 = {1{`RANDOM}};
  lineBuffer_674 = _RAND_681[7:0];
  _RAND_682 = {1{`RANDOM}};
  lineBuffer_675 = _RAND_682[7:0];
  _RAND_683 = {1{`RANDOM}};
  lineBuffer_676 = _RAND_683[7:0];
  _RAND_684 = {1{`RANDOM}};
  lineBuffer_677 = _RAND_684[7:0];
  _RAND_685 = {1{`RANDOM}};
  lineBuffer_678 = _RAND_685[7:0];
  _RAND_686 = {1{`RANDOM}};
  lineBuffer_679 = _RAND_686[7:0];
  _RAND_687 = {1{`RANDOM}};
  lineBuffer_680 = _RAND_687[7:0];
  _RAND_688 = {1{`RANDOM}};
  lineBuffer_681 = _RAND_688[7:0];
  _RAND_689 = {1{`RANDOM}};
  lineBuffer_682 = _RAND_689[7:0];
  _RAND_690 = {1{`RANDOM}};
  lineBuffer_683 = _RAND_690[7:0];
  _RAND_691 = {1{`RANDOM}};
  lineBuffer_684 = _RAND_691[7:0];
  _RAND_692 = {1{`RANDOM}};
  lineBuffer_685 = _RAND_692[7:0];
  _RAND_693 = {1{`RANDOM}};
  lineBuffer_686 = _RAND_693[7:0];
  _RAND_694 = {1{`RANDOM}};
  lineBuffer_687 = _RAND_694[7:0];
  _RAND_695 = {1{`RANDOM}};
  lineBuffer_688 = _RAND_695[7:0];
  _RAND_696 = {1{`RANDOM}};
  lineBuffer_689 = _RAND_696[7:0];
  _RAND_697 = {1{`RANDOM}};
  lineBuffer_690 = _RAND_697[7:0];
  _RAND_698 = {1{`RANDOM}};
  lineBuffer_691 = _RAND_698[7:0];
  _RAND_699 = {1{`RANDOM}};
  lineBuffer_692 = _RAND_699[7:0];
  _RAND_700 = {1{`RANDOM}};
  lineBuffer_693 = _RAND_700[7:0];
  _RAND_701 = {1{`RANDOM}};
  lineBuffer_694 = _RAND_701[7:0];
  _RAND_702 = {1{`RANDOM}};
  lineBuffer_695 = _RAND_702[7:0];
  _RAND_703 = {1{`RANDOM}};
  lineBuffer_696 = _RAND_703[7:0];
  _RAND_704 = {1{`RANDOM}};
  lineBuffer_697 = _RAND_704[7:0];
  _RAND_705 = {1{`RANDOM}};
  lineBuffer_698 = _RAND_705[7:0];
  _RAND_706 = {1{`RANDOM}};
  lineBuffer_699 = _RAND_706[7:0];
  _RAND_707 = {1{`RANDOM}};
  lineBuffer_700 = _RAND_707[7:0];
  _RAND_708 = {1{`RANDOM}};
  lineBuffer_701 = _RAND_708[7:0];
  _RAND_709 = {1{`RANDOM}};
  lineBuffer_702 = _RAND_709[7:0];
  _RAND_710 = {1{`RANDOM}};
  lineBuffer_703 = _RAND_710[7:0];
  _RAND_711 = {1{`RANDOM}};
  lineBuffer_704 = _RAND_711[7:0];
  _RAND_712 = {1{`RANDOM}};
  lineBuffer_705 = _RAND_712[7:0];
  _RAND_713 = {1{`RANDOM}};
  lineBuffer_706 = _RAND_713[7:0];
  _RAND_714 = {1{`RANDOM}};
  lineBuffer_707 = _RAND_714[7:0];
  _RAND_715 = {1{`RANDOM}};
  lineBuffer_708 = _RAND_715[7:0];
  _RAND_716 = {1{`RANDOM}};
  lineBuffer_709 = _RAND_716[7:0];
  _RAND_717 = {1{`RANDOM}};
  lineBuffer_710 = _RAND_717[7:0];
  _RAND_718 = {1{`RANDOM}};
  lineBuffer_711 = _RAND_718[7:0];
  _RAND_719 = {1{`RANDOM}};
  lineBuffer_712 = _RAND_719[7:0];
  _RAND_720 = {1{`RANDOM}};
  lineBuffer_713 = _RAND_720[7:0];
  _RAND_721 = {1{`RANDOM}};
  lineBuffer_714 = _RAND_721[7:0];
  _RAND_722 = {1{`RANDOM}};
  lineBuffer_715 = _RAND_722[7:0];
  _RAND_723 = {1{`RANDOM}};
  lineBuffer_716 = _RAND_723[7:0];
  _RAND_724 = {1{`RANDOM}};
  lineBuffer_717 = _RAND_724[7:0];
  _RAND_725 = {1{`RANDOM}};
  lineBuffer_718 = _RAND_725[7:0];
  _RAND_726 = {1{`RANDOM}};
  lineBuffer_719 = _RAND_726[7:0];
  _RAND_727 = {1{`RANDOM}};
  lineBuffer_720 = _RAND_727[7:0];
  _RAND_728 = {1{`RANDOM}};
  lineBuffer_721 = _RAND_728[7:0];
  _RAND_729 = {1{`RANDOM}};
  lineBuffer_722 = _RAND_729[7:0];
  _RAND_730 = {1{`RANDOM}};
  lineBuffer_723 = _RAND_730[7:0];
  _RAND_731 = {1{`RANDOM}};
  lineBuffer_724 = _RAND_731[7:0];
  _RAND_732 = {1{`RANDOM}};
  lineBuffer_725 = _RAND_732[7:0];
  _RAND_733 = {1{`RANDOM}};
  lineBuffer_726 = _RAND_733[7:0];
  _RAND_734 = {1{`RANDOM}};
  lineBuffer_727 = _RAND_734[7:0];
  _RAND_735 = {1{`RANDOM}};
  lineBuffer_728 = _RAND_735[7:0];
  _RAND_736 = {1{`RANDOM}};
  lineBuffer_729 = _RAND_736[7:0];
  _RAND_737 = {1{`RANDOM}};
  lineBuffer_730 = _RAND_737[7:0];
  _RAND_738 = {1{`RANDOM}};
  lineBuffer_731 = _RAND_738[7:0];
  _RAND_739 = {1{`RANDOM}};
  lineBuffer_732 = _RAND_739[7:0];
  _RAND_740 = {1{`RANDOM}};
  lineBuffer_733 = _RAND_740[7:0];
  _RAND_741 = {1{`RANDOM}};
  lineBuffer_734 = _RAND_741[7:0];
  _RAND_742 = {1{`RANDOM}};
  lineBuffer_735 = _RAND_742[7:0];
  _RAND_743 = {1{`RANDOM}};
  lineBuffer_736 = _RAND_743[7:0];
  _RAND_744 = {1{`RANDOM}};
  lineBuffer_737 = _RAND_744[7:0];
  _RAND_745 = {1{`RANDOM}};
  lineBuffer_738 = _RAND_745[7:0];
  _RAND_746 = {1{`RANDOM}};
  lineBuffer_739 = _RAND_746[7:0];
  _RAND_747 = {1{`RANDOM}};
  lineBuffer_740 = _RAND_747[7:0];
  _RAND_748 = {1{`RANDOM}};
  lineBuffer_741 = _RAND_748[7:0];
  _RAND_749 = {1{`RANDOM}};
  lineBuffer_742 = _RAND_749[7:0];
  _RAND_750 = {1{`RANDOM}};
  lineBuffer_743 = _RAND_750[7:0];
  _RAND_751 = {1{`RANDOM}};
  lineBuffer_744 = _RAND_751[7:0];
  _RAND_752 = {1{`RANDOM}};
  lineBuffer_745 = _RAND_752[7:0];
  _RAND_753 = {1{`RANDOM}};
  lineBuffer_746 = _RAND_753[7:0];
  _RAND_754 = {1{`RANDOM}};
  lineBuffer_747 = _RAND_754[7:0];
  _RAND_755 = {1{`RANDOM}};
  lineBuffer_748 = _RAND_755[7:0];
  _RAND_756 = {1{`RANDOM}};
  lineBuffer_749 = _RAND_756[7:0];
  _RAND_757 = {1{`RANDOM}};
  lineBuffer_750 = _RAND_757[7:0];
  _RAND_758 = {1{`RANDOM}};
  lineBuffer_751 = _RAND_758[7:0];
  _RAND_759 = {1{`RANDOM}};
  lineBuffer_752 = _RAND_759[7:0];
  _RAND_760 = {1{`RANDOM}};
  lineBuffer_753 = _RAND_760[7:0];
  _RAND_761 = {1{`RANDOM}};
  lineBuffer_754 = _RAND_761[7:0];
  _RAND_762 = {1{`RANDOM}};
  lineBuffer_755 = _RAND_762[7:0];
  _RAND_763 = {1{`RANDOM}};
  lineBuffer_756 = _RAND_763[7:0];
  _RAND_764 = {1{`RANDOM}};
  lineBuffer_757 = _RAND_764[7:0];
  _RAND_765 = {1{`RANDOM}};
  lineBuffer_758 = _RAND_765[7:0];
  _RAND_766 = {1{`RANDOM}};
  lineBuffer_759 = _RAND_766[7:0];
  _RAND_767 = {1{`RANDOM}};
  lineBuffer_760 = _RAND_767[7:0];
  _RAND_768 = {1{`RANDOM}};
  lineBuffer_761 = _RAND_768[7:0];
  _RAND_769 = {1{`RANDOM}};
  lineBuffer_762 = _RAND_769[7:0];
  _RAND_770 = {1{`RANDOM}};
  lineBuffer_763 = _RAND_770[7:0];
  _RAND_771 = {1{`RANDOM}};
  lineBuffer_764 = _RAND_771[7:0];
  _RAND_772 = {1{`RANDOM}};
  lineBuffer_765 = _RAND_772[7:0];
  _RAND_773 = {1{`RANDOM}};
  lineBuffer_766 = _RAND_773[7:0];
  _RAND_774 = {1{`RANDOM}};
  lineBuffer_767 = _RAND_774[7:0];
  _RAND_775 = {1{`RANDOM}};
  windowBuffer_0 = _RAND_775[7:0];
  _RAND_776 = {1{`RANDOM}};
  windowBuffer_1 = _RAND_776[7:0];
  _RAND_777 = {1{`RANDOM}};
  windowBuffer_2 = _RAND_777[7:0];
  _RAND_778 = {1{`RANDOM}};
  windowBuffer_3 = _RAND_778[7:0];
  _RAND_779 = {1{`RANDOM}};
  windowBuffer_4 = _RAND_779[7:0];
  _RAND_780 = {1{`RANDOM}};
  windowBuffer_5 = _RAND_780[7:0];
  _RAND_781 = {1{`RANDOM}};
  windowBuffer_6 = _RAND_781[7:0];
  _RAND_782 = {1{`RANDOM}};
  windowBuffer_7 = _RAND_782[7:0];
  _RAND_783 = {1{`RANDOM}};
  windowBuffer_8 = _RAND_783[7:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      stateReg <= 2'h0;
    end else if (_T) begin
      if (io__enq_valid) begin
        stateReg <= 2'h1;
      end
    end else if (_T_1) begin
      if (_T_3) begin
        stateReg <= 2'h0;
      end else if (_T_4) begin
        stateReg <= 2'h1;
      end else if (_T_6) begin
        stateReg <= 2'h2;
      end
    end else if (_T_7) begin
      if (io__deq_ready) begin
        stateReg <= 2'h1;
      end
    end else if (_T_8) begin
      stateReg <= 2'h0;
    end
    if (_T) begin
      if (io__enq_valid) begin
        dataReg <= io__enq_bits;
      end
    end else if (_T_1) begin
      if (!(_T_3)) begin
        if (_T_4) begin
          dataReg <= io__enq_bits;
        end
      end
    end else if (_T_7) begin
      if (io__deq_ready) begin
        dataReg <= shadowReg;
      end
    end
    if (!(_T)) begin
      if (_T_1) begin
        if (!(_T_3)) begin
          if (!(_T_4)) begin
            if (_T_6) begin
              shadowReg <= io__enq_bits;
            end
          end
        end
      end
    end
    if (_T) begin
      userReg <= io__enq_user;
    end else if (_T_1) begin
      if (_T_3) begin
        userReg <= io__enq_user;
      end else if (_T_4) begin
        userReg <= io__enq_user;
      end
    end else if (_T_7) begin
      if (io__deq_ready) begin
        userReg <= shadowUserReg;
      end
    end
    if (!(_T)) begin
      if (_T_1) begin
        if (!(_T_3)) begin
          if (!(_T_4)) begin
            if (_T_6) begin
              shadowUserReg <= io__enq_user;
            end
          end
        end
      end
    end
    if (_T) begin
      if (io__enq_valid) begin
        lastReg <= io__enq_last;
      end
    end else if (_T_1) begin
      if (!(_T_3)) begin
        if (_T_4) begin
          lastReg <= io__enq_last;
        end
      end
    end else if (_T_7) begin
      if (io__deq_ready) begin
        lastReg <= shadowLastReg;
      end
    end
    if (!(_T)) begin
      if (_T_1) begin
        if (!(_T_3)) begin
          if (!(_T_4)) begin
            if (_T_6) begin
              shadowLastReg <= io__enq_last;
            end
          end
        end
      end
    end
    if (sel) begin
      lineBuffer_0 <= dataReg;
    end
    if (sel) begin
      lineBuffer_1 <= lineBuffer_0;
    end
    if (sel) begin
      lineBuffer_2 <= lineBuffer_1;
    end
    if (sel) begin
      lineBuffer_3 <= lineBuffer_2;
    end
    if (sel) begin
      lineBuffer_4 <= lineBuffer_3;
    end
    if (sel) begin
      lineBuffer_5 <= lineBuffer_4;
    end
    if (sel) begin
      lineBuffer_6 <= lineBuffer_5;
    end
    if (sel) begin
      lineBuffer_7 <= lineBuffer_6;
    end
    if (sel) begin
      lineBuffer_8 <= lineBuffer_7;
    end
    if (sel) begin
      lineBuffer_9 <= lineBuffer_8;
    end
    if (sel) begin
      lineBuffer_10 <= lineBuffer_9;
    end
    if (sel) begin
      lineBuffer_11 <= lineBuffer_10;
    end
    if (sel) begin
      lineBuffer_12 <= lineBuffer_11;
    end
    if (sel) begin
      lineBuffer_13 <= lineBuffer_12;
    end
    if (sel) begin
      lineBuffer_14 <= lineBuffer_13;
    end
    if (sel) begin
      lineBuffer_15 <= lineBuffer_14;
    end
    if (sel) begin
      lineBuffer_16 <= lineBuffer_15;
    end
    if (sel) begin
      lineBuffer_17 <= lineBuffer_16;
    end
    if (sel) begin
      lineBuffer_18 <= lineBuffer_17;
    end
    if (sel) begin
      lineBuffer_19 <= lineBuffer_18;
    end
    if (sel) begin
      lineBuffer_20 <= lineBuffer_19;
    end
    if (sel) begin
      lineBuffer_21 <= lineBuffer_20;
    end
    if (sel) begin
      lineBuffer_22 <= lineBuffer_21;
    end
    if (sel) begin
      lineBuffer_23 <= lineBuffer_22;
    end
    if (sel) begin
      lineBuffer_24 <= lineBuffer_23;
    end
    if (sel) begin
      lineBuffer_25 <= lineBuffer_24;
    end
    if (sel) begin
      lineBuffer_26 <= lineBuffer_25;
    end
    if (sel) begin
      lineBuffer_27 <= lineBuffer_26;
    end
    if (sel) begin
      lineBuffer_28 <= lineBuffer_27;
    end
    if (sel) begin
      lineBuffer_29 <= lineBuffer_28;
    end
    if (sel) begin
      lineBuffer_30 <= lineBuffer_29;
    end
    if (sel) begin
      lineBuffer_31 <= lineBuffer_30;
    end
    if (sel) begin
      lineBuffer_32 <= lineBuffer_31;
    end
    if (sel) begin
      lineBuffer_33 <= lineBuffer_32;
    end
    if (sel) begin
      lineBuffer_34 <= lineBuffer_33;
    end
    if (sel) begin
      lineBuffer_35 <= lineBuffer_34;
    end
    if (sel) begin
      lineBuffer_36 <= lineBuffer_35;
    end
    if (sel) begin
      lineBuffer_37 <= lineBuffer_36;
    end
    if (sel) begin
      lineBuffer_38 <= lineBuffer_37;
    end
    if (sel) begin
      lineBuffer_39 <= lineBuffer_38;
    end
    if (sel) begin
      lineBuffer_40 <= lineBuffer_39;
    end
    if (sel) begin
      lineBuffer_41 <= lineBuffer_40;
    end
    if (sel) begin
      lineBuffer_42 <= lineBuffer_41;
    end
    if (sel) begin
      lineBuffer_43 <= lineBuffer_42;
    end
    if (sel) begin
      lineBuffer_44 <= lineBuffer_43;
    end
    if (sel) begin
      lineBuffer_45 <= lineBuffer_44;
    end
    if (sel) begin
      lineBuffer_46 <= lineBuffer_45;
    end
    if (sel) begin
      lineBuffer_47 <= lineBuffer_46;
    end
    if (sel) begin
      lineBuffer_48 <= lineBuffer_47;
    end
    if (sel) begin
      lineBuffer_49 <= lineBuffer_48;
    end
    if (sel) begin
      lineBuffer_50 <= lineBuffer_49;
    end
    if (sel) begin
      lineBuffer_51 <= lineBuffer_50;
    end
    if (sel) begin
      lineBuffer_52 <= lineBuffer_51;
    end
    if (sel) begin
      lineBuffer_53 <= lineBuffer_52;
    end
    if (sel) begin
      lineBuffer_54 <= lineBuffer_53;
    end
    if (sel) begin
      lineBuffer_55 <= lineBuffer_54;
    end
    if (sel) begin
      lineBuffer_56 <= lineBuffer_55;
    end
    if (sel) begin
      lineBuffer_57 <= lineBuffer_56;
    end
    if (sel) begin
      lineBuffer_58 <= lineBuffer_57;
    end
    if (sel) begin
      lineBuffer_59 <= lineBuffer_58;
    end
    if (sel) begin
      lineBuffer_60 <= lineBuffer_59;
    end
    if (sel) begin
      lineBuffer_61 <= lineBuffer_60;
    end
    if (sel) begin
      lineBuffer_62 <= lineBuffer_61;
    end
    if (sel) begin
      lineBuffer_63 <= lineBuffer_62;
    end
    if (sel) begin
      lineBuffer_64 <= lineBuffer_63;
    end
    if (sel) begin
      lineBuffer_65 <= lineBuffer_64;
    end
    if (sel) begin
      lineBuffer_66 <= lineBuffer_65;
    end
    if (sel) begin
      lineBuffer_67 <= lineBuffer_66;
    end
    if (sel) begin
      lineBuffer_68 <= lineBuffer_67;
    end
    if (sel) begin
      lineBuffer_69 <= lineBuffer_68;
    end
    if (sel) begin
      lineBuffer_70 <= lineBuffer_69;
    end
    if (sel) begin
      lineBuffer_71 <= lineBuffer_70;
    end
    if (sel) begin
      lineBuffer_72 <= lineBuffer_71;
    end
    if (sel) begin
      lineBuffer_73 <= lineBuffer_72;
    end
    if (sel) begin
      lineBuffer_74 <= lineBuffer_73;
    end
    if (sel) begin
      lineBuffer_75 <= lineBuffer_74;
    end
    if (sel) begin
      lineBuffer_76 <= lineBuffer_75;
    end
    if (sel) begin
      lineBuffer_77 <= lineBuffer_76;
    end
    if (sel) begin
      lineBuffer_78 <= lineBuffer_77;
    end
    if (sel) begin
      lineBuffer_79 <= lineBuffer_78;
    end
    if (sel) begin
      lineBuffer_80 <= lineBuffer_79;
    end
    if (sel) begin
      lineBuffer_81 <= lineBuffer_80;
    end
    if (sel) begin
      lineBuffer_82 <= lineBuffer_81;
    end
    if (sel) begin
      lineBuffer_83 <= lineBuffer_82;
    end
    if (sel) begin
      lineBuffer_84 <= lineBuffer_83;
    end
    if (sel) begin
      lineBuffer_85 <= lineBuffer_84;
    end
    if (sel) begin
      lineBuffer_86 <= lineBuffer_85;
    end
    if (sel) begin
      lineBuffer_87 <= lineBuffer_86;
    end
    if (sel) begin
      lineBuffer_88 <= lineBuffer_87;
    end
    if (sel) begin
      lineBuffer_89 <= lineBuffer_88;
    end
    if (sel) begin
      lineBuffer_90 <= lineBuffer_89;
    end
    if (sel) begin
      lineBuffer_91 <= lineBuffer_90;
    end
    if (sel) begin
      lineBuffer_92 <= lineBuffer_91;
    end
    if (sel) begin
      lineBuffer_93 <= lineBuffer_92;
    end
    if (sel) begin
      lineBuffer_94 <= lineBuffer_93;
    end
    if (sel) begin
      lineBuffer_95 <= lineBuffer_94;
    end
    if (sel) begin
      lineBuffer_96 <= lineBuffer_95;
    end
    if (sel) begin
      lineBuffer_97 <= lineBuffer_96;
    end
    if (sel) begin
      lineBuffer_98 <= lineBuffer_97;
    end
    if (sel) begin
      lineBuffer_99 <= lineBuffer_98;
    end
    if (sel) begin
      lineBuffer_100 <= lineBuffer_99;
    end
    if (sel) begin
      lineBuffer_101 <= lineBuffer_100;
    end
    if (sel) begin
      lineBuffer_102 <= lineBuffer_101;
    end
    if (sel) begin
      lineBuffer_103 <= lineBuffer_102;
    end
    if (sel) begin
      lineBuffer_104 <= lineBuffer_103;
    end
    if (sel) begin
      lineBuffer_105 <= lineBuffer_104;
    end
    if (sel) begin
      lineBuffer_106 <= lineBuffer_105;
    end
    if (sel) begin
      lineBuffer_107 <= lineBuffer_106;
    end
    if (sel) begin
      lineBuffer_108 <= lineBuffer_107;
    end
    if (sel) begin
      lineBuffer_109 <= lineBuffer_108;
    end
    if (sel) begin
      lineBuffer_110 <= lineBuffer_109;
    end
    if (sel) begin
      lineBuffer_111 <= lineBuffer_110;
    end
    if (sel) begin
      lineBuffer_112 <= lineBuffer_111;
    end
    if (sel) begin
      lineBuffer_113 <= lineBuffer_112;
    end
    if (sel) begin
      lineBuffer_114 <= lineBuffer_113;
    end
    if (sel) begin
      lineBuffer_115 <= lineBuffer_114;
    end
    if (sel) begin
      lineBuffer_116 <= lineBuffer_115;
    end
    if (sel) begin
      lineBuffer_117 <= lineBuffer_116;
    end
    if (sel) begin
      lineBuffer_118 <= lineBuffer_117;
    end
    if (sel) begin
      lineBuffer_119 <= lineBuffer_118;
    end
    if (sel) begin
      lineBuffer_120 <= lineBuffer_119;
    end
    if (sel) begin
      lineBuffer_121 <= lineBuffer_120;
    end
    if (sel) begin
      lineBuffer_122 <= lineBuffer_121;
    end
    if (sel) begin
      lineBuffer_123 <= lineBuffer_122;
    end
    if (sel) begin
      lineBuffer_124 <= lineBuffer_123;
    end
    if (sel) begin
      lineBuffer_125 <= lineBuffer_124;
    end
    if (sel) begin
      lineBuffer_126 <= lineBuffer_125;
    end
    if (sel) begin
      lineBuffer_127 <= lineBuffer_126;
    end
    if (sel) begin
      lineBuffer_128 <= lineBuffer_127;
    end
    if (sel) begin
      lineBuffer_129 <= lineBuffer_128;
    end
    if (sel) begin
      lineBuffer_130 <= lineBuffer_129;
    end
    if (sel) begin
      lineBuffer_131 <= lineBuffer_130;
    end
    if (sel) begin
      lineBuffer_132 <= lineBuffer_131;
    end
    if (sel) begin
      lineBuffer_133 <= lineBuffer_132;
    end
    if (sel) begin
      lineBuffer_134 <= lineBuffer_133;
    end
    if (sel) begin
      lineBuffer_135 <= lineBuffer_134;
    end
    if (sel) begin
      lineBuffer_136 <= lineBuffer_135;
    end
    if (sel) begin
      lineBuffer_137 <= lineBuffer_136;
    end
    if (sel) begin
      lineBuffer_138 <= lineBuffer_137;
    end
    if (sel) begin
      lineBuffer_139 <= lineBuffer_138;
    end
    if (sel) begin
      lineBuffer_140 <= lineBuffer_139;
    end
    if (sel) begin
      lineBuffer_141 <= lineBuffer_140;
    end
    if (sel) begin
      lineBuffer_142 <= lineBuffer_141;
    end
    if (sel) begin
      lineBuffer_143 <= lineBuffer_142;
    end
    if (sel) begin
      lineBuffer_144 <= lineBuffer_143;
    end
    if (sel) begin
      lineBuffer_145 <= lineBuffer_144;
    end
    if (sel) begin
      lineBuffer_146 <= lineBuffer_145;
    end
    if (sel) begin
      lineBuffer_147 <= lineBuffer_146;
    end
    if (sel) begin
      lineBuffer_148 <= lineBuffer_147;
    end
    if (sel) begin
      lineBuffer_149 <= lineBuffer_148;
    end
    if (sel) begin
      lineBuffer_150 <= lineBuffer_149;
    end
    if (sel) begin
      lineBuffer_151 <= lineBuffer_150;
    end
    if (sel) begin
      lineBuffer_152 <= lineBuffer_151;
    end
    if (sel) begin
      lineBuffer_153 <= lineBuffer_152;
    end
    if (sel) begin
      lineBuffer_154 <= lineBuffer_153;
    end
    if (sel) begin
      lineBuffer_155 <= lineBuffer_154;
    end
    if (sel) begin
      lineBuffer_156 <= lineBuffer_155;
    end
    if (sel) begin
      lineBuffer_157 <= lineBuffer_156;
    end
    if (sel) begin
      lineBuffer_158 <= lineBuffer_157;
    end
    if (sel) begin
      lineBuffer_159 <= lineBuffer_158;
    end
    if (sel) begin
      lineBuffer_160 <= lineBuffer_159;
    end
    if (sel) begin
      lineBuffer_161 <= lineBuffer_160;
    end
    if (sel) begin
      lineBuffer_162 <= lineBuffer_161;
    end
    if (sel) begin
      lineBuffer_163 <= lineBuffer_162;
    end
    if (sel) begin
      lineBuffer_164 <= lineBuffer_163;
    end
    if (sel) begin
      lineBuffer_165 <= lineBuffer_164;
    end
    if (sel) begin
      lineBuffer_166 <= lineBuffer_165;
    end
    if (sel) begin
      lineBuffer_167 <= lineBuffer_166;
    end
    if (sel) begin
      lineBuffer_168 <= lineBuffer_167;
    end
    if (sel) begin
      lineBuffer_169 <= lineBuffer_168;
    end
    if (sel) begin
      lineBuffer_170 <= lineBuffer_169;
    end
    if (sel) begin
      lineBuffer_171 <= lineBuffer_170;
    end
    if (sel) begin
      lineBuffer_172 <= lineBuffer_171;
    end
    if (sel) begin
      lineBuffer_173 <= lineBuffer_172;
    end
    if (sel) begin
      lineBuffer_174 <= lineBuffer_173;
    end
    if (sel) begin
      lineBuffer_175 <= lineBuffer_174;
    end
    if (sel) begin
      lineBuffer_176 <= lineBuffer_175;
    end
    if (sel) begin
      lineBuffer_177 <= lineBuffer_176;
    end
    if (sel) begin
      lineBuffer_178 <= lineBuffer_177;
    end
    if (sel) begin
      lineBuffer_179 <= lineBuffer_178;
    end
    if (sel) begin
      lineBuffer_180 <= lineBuffer_179;
    end
    if (sel) begin
      lineBuffer_181 <= lineBuffer_180;
    end
    if (sel) begin
      lineBuffer_182 <= lineBuffer_181;
    end
    if (sel) begin
      lineBuffer_183 <= lineBuffer_182;
    end
    if (sel) begin
      lineBuffer_184 <= lineBuffer_183;
    end
    if (sel) begin
      lineBuffer_185 <= lineBuffer_184;
    end
    if (sel) begin
      lineBuffer_186 <= lineBuffer_185;
    end
    if (sel) begin
      lineBuffer_187 <= lineBuffer_186;
    end
    if (sel) begin
      lineBuffer_188 <= lineBuffer_187;
    end
    if (sel) begin
      lineBuffer_189 <= lineBuffer_188;
    end
    if (sel) begin
      lineBuffer_190 <= lineBuffer_189;
    end
    if (sel) begin
      lineBuffer_191 <= lineBuffer_190;
    end
    if (sel) begin
      lineBuffer_192 <= lineBuffer_191;
    end
    if (sel) begin
      lineBuffer_193 <= lineBuffer_192;
    end
    if (sel) begin
      lineBuffer_194 <= lineBuffer_193;
    end
    if (sel) begin
      lineBuffer_195 <= lineBuffer_194;
    end
    if (sel) begin
      lineBuffer_196 <= lineBuffer_195;
    end
    if (sel) begin
      lineBuffer_197 <= lineBuffer_196;
    end
    if (sel) begin
      lineBuffer_198 <= lineBuffer_197;
    end
    if (sel) begin
      lineBuffer_199 <= lineBuffer_198;
    end
    if (sel) begin
      lineBuffer_200 <= lineBuffer_199;
    end
    if (sel) begin
      lineBuffer_201 <= lineBuffer_200;
    end
    if (sel) begin
      lineBuffer_202 <= lineBuffer_201;
    end
    if (sel) begin
      lineBuffer_203 <= lineBuffer_202;
    end
    if (sel) begin
      lineBuffer_204 <= lineBuffer_203;
    end
    if (sel) begin
      lineBuffer_205 <= lineBuffer_204;
    end
    if (sel) begin
      lineBuffer_206 <= lineBuffer_205;
    end
    if (sel) begin
      lineBuffer_207 <= lineBuffer_206;
    end
    if (sel) begin
      lineBuffer_208 <= lineBuffer_207;
    end
    if (sel) begin
      lineBuffer_209 <= lineBuffer_208;
    end
    if (sel) begin
      lineBuffer_210 <= lineBuffer_209;
    end
    if (sel) begin
      lineBuffer_211 <= lineBuffer_210;
    end
    if (sel) begin
      lineBuffer_212 <= lineBuffer_211;
    end
    if (sel) begin
      lineBuffer_213 <= lineBuffer_212;
    end
    if (sel) begin
      lineBuffer_214 <= lineBuffer_213;
    end
    if (sel) begin
      lineBuffer_215 <= lineBuffer_214;
    end
    if (sel) begin
      lineBuffer_216 <= lineBuffer_215;
    end
    if (sel) begin
      lineBuffer_217 <= lineBuffer_216;
    end
    if (sel) begin
      lineBuffer_218 <= lineBuffer_217;
    end
    if (sel) begin
      lineBuffer_219 <= lineBuffer_218;
    end
    if (sel) begin
      lineBuffer_220 <= lineBuffer_219;
    end
    if (sel) begin
      lineBuffer_221 <= lineBuffer_220;
    end
    if (sel) begin
      lineBuffer_222 <= lineBuffer_221;
    end
    if (sel) begin
      lineBuffer_223 <= lineBuffer_222;
    end
    if (sel) begin
      lineBuffer_224 <= lineBuffer_223;
    end
    if (sel) begin
      lineBuffer_225 <= lineBuffer_224;
    end
    if (sel) begin
      lineBuffer_226 <= lineBuffer_225;
    end
    if (sel) begin
      lineBuffer_227 <= lineBuffer_226;
    end
    if (sel) begin
      lineBuffer_228 <= lineBuffer_227;
    end
    if (sel) begin
      lineBuffer_229 <= lineBuffer_228;
    end
    if (sel) begin
      lineBuffer_230 <= lineBuffer_229;
    end
    if (sel) begin
      lineBuffer_231 <= lineBuffer_230;
    end
    if (sel) begin
      lineBuffer_232 <= lineBuffer_231;
    end
    if (sel) begin
      lineBuffer_233 <= lineBuffer_232;
    end
    if (sel) begin
      lineBuffer_234 <= lineBuffer_233;
    end
    if (sel) begin
      lineBuffer_235 <= lineBuffer_234;
    end
    if (sel) begin
      lineBuffer_236 <= lineBuffer_235;
    end
    if (sel) begin
      lineBuffer_237 <= lineBuffer_236;
    end
    if (sel) begin
      lineBuffer_238 <= lineBuffer_237;
    end
    if (sel) begin
      lineBuffer_239 <= lineBuffer_238;
    end
    if (sel) begin
      lineBuffer_240 <= lineBuffer_239;
    end
    if (sel) begin
      lineBuffer_241 <= lineBuffer_240;
    end
    if (sel) begin
      lineBuffer_242 <= lineBuffer_241;
    end
    if (sel) begin
      lineBuffer_243 <= lineBuffer_242;
    end
    if (sel) begin
      lineBuffer_244 <= lineBuffer_243;
    end
    if (sel) begin
      lineBuffer_245 <= lineBuffer_244;
    end
    if (sel) begin
      lineBuffer_246 <= lineBuffer_245;
    end
    if (sel) begin
      lineBuffer_247 <= lineBuffer_246;
    end
    if (sel) begin
      lineBuffer_248 <= lineBuffer_247;
    end
    if (sel) begin
      lineBuffer_249 <= lineBuffer_248;
    end
    if (sel) begin
      lineBuffer_250 <= lineBuffer_249;
    end
    if (sel) begin
      lineBuffer_251 <= lineBuffer_250;
    end
    if (sel) begin
      lineBuffer_252 <= lineBuffer_251;
    end
    if (sel) begin
      lineBuffer_253 <= lineBuffer_252;
    end
    if (sel) begin
      lineBuffer_254 <= lineBuffer_253;
    end
    if (sel) begin
      lineBuffer_255 <= lineBuffer_254;
    end
    if (sel) begin
      lineBuffer_256 <= lineBuffer_255;
    end
    if (sel) begin
      lineBuffer_257 <= lineBuffer_256;
    end
    if (sel) begin
      lineBuffer_258 <= lineBuffer_257;
    end
    if (sel) begin
      lineBuffer_259 <= lineBuffer_258;
    end
    if (sel) begin
      lineBuffer_260 <= lineBuffer_259;
    end
    if (sel) begin
      lineBuffer_261 <= lineBuffer_260;
    end
    if (sel) begin
      lineBuffer_262 <= lineBuffer_261;
    end
    if (sel) begin
      lineBuffer_263 <= lineBuffer_262;
    end
    if (sel) begin
      lineBuffer_264 <= lineBuffer_263;
    end
    if (sel) begin
      lineBuffer_265 <= lineBuffer_264;
    end
    if (sel) begin
      lineBuffer_266 <= lineBuffer_265;
    end
    if (sel) begin
      lineBuffer_267 <= lineBuffer_266;
    end
    if (sel) begin
      lineBuffer_268 <= lineBuffer_267;
    end
    if (sel) begin
      lineBuffer_269 <= lineBuffer_268;
    end
    if (sel) begin
      lineBuffer_270 <= lineBuffer_269;
    end
    if (sel) begin
      lineBuffer_271 <= lineBuffer_270;
    end
    if (sel) begin
      lineBuffer_272 <= lineBuffer_271;
    end
    if (sel) begin
      lineBuffer_273 <= lineBuffer_272;
    end
    if (sel) begin
      lineBuffer_274 <= lineBuffer_273;
    end
    if (sel) begin
      lineBuffer_275 <= lineBuffer_274;
    end
    if (sel) begin
      lineBuffer_276 <= lineBuffer_275;
    end
    if (sel) begin
      lineBuffer_277 <= lineBuffer_276;
    end
    if (sel) begin
      lineBuffer_278 <= lineBuffer_277;
    end
    if (sel) begin
      lineBuffer_279 <= lineBuffer_278;
    end
    if (sel) begin
      lineBuffer_280 <= lineBuffer_279;
    end
    if (sel) begin
      lineBuffer_281 <= lineBuffer_280;
    end
    if (sel) begin
      lineBuffer_282 <= lineBuffer_281;
    end
    if (sel) begin
      lineBuffer_283 <= lineBuffer_282;
    end
    if (sel) begin
      lineBuffer_284 <= lineBuffer_283;
    end
    if (sel) begin
      lineBuffer_285 <= lineBuffer_284;
    end
    if (sel) begin
      lineBuffer_286 <= lineBuffer_285;
    end
    if (sel) begin
      lineBuffer_287 <= lineBuffer_286;
    end
    if (sel) begin
      lineBuffer_288 <= lineBuffer_287;
    end
    if (sel) begin
      lineBuffer_289 <= lineBuffer_288;
    end
    if (sel) begin
      lineBuffer_290 <= lineBuffer_289;
    end
    if (sel) begin
      lineBuffer_291 <= lineBuffer_290;
    end
    if (sel) begin
      lineBuffer_292 <= lineBuffer_291;
    end
    if (sel) begin
      lineBuffer_293 <= lineBuffer_292;
    end
    if (sel) begin
      lineBuffer_294 <= lineBuffer_293;
    end
    if (sel) begin
      lineBuffer_295 <= lineBuffer_294;
    end
    if (sel) begin
      lineBuffer_296 <= lineBuffer_295;
    end
    if (sel) begin
      lineBuffer_297 <= lineBuffer_296;
    end
    if (sel) begin
      lineBuffer_298 <= lineBuffer_297;
    end
    if (sel) begin
      lineBuffer_299 <= lineBuffer_298;
    end
    if (sel) begin
      lineBuffer_300 <= lineBuffer_299;
    end
    if (sel) begin
      lineBuffer_301 <= lineBuffer_300;
    end
    if (sel) begin
      lineBuffer_302 <= lineBuffer_301;
    end
    if (sel) begin
      lineBuffer_303 <= lineBuffer_302;
    end
    if (sel) begin
      lineBuffer_304 <= lineBuffer_303;
    end
    if (sel) begin
      lineBuffer_305 <= lineBuffer_304;
    end
    if (sel) begin
      lineBuffer_306 <= lineBuffer_305;
    end
    if (sel) begin
      lineBuffer_307 <= lineBuffer_306;
    end
    if (sel) begin
      lineBuffer_308 <= lineBuffer_307;
    end
    if (sel) begin
      lineBuffer_309 <= lineBuffer_308;
    end
    if (sel) begin
      lineBuffer_310 <= lineBuffer_309;
    end
    if (sel) begin
      lineBuffer_311 <= lineBuffer_310;
    end
    if (sel) begin
      lineBuffer_312 <= lineBuffer_311;
    end
    if (sel) begin
      lineBuffer_313 <= lineBuffer_312;
    end
    if (sel) begin
      lineBuffer_314 <= lineBuffer_313;
    end
    if (sel) begin
      lineBuffer_315 <= lineBuffer_314;
    end
    if (sel) begin
      lineBuffer_316 <= lineBuffer_315;
    end
    if (sel) begin
      lineBuffer_317 <= lineBuffer_316;
    end
    if (sel) begin
      lineBuffer_318 <= lineBuffer_317;
    end
    if (sel) begin
      lineBuffer_319 <= lineBuffer_318;
    end
    if (sel) begin
      lineBuffer_320 <= lineBuffer_319;
    end
    if (sel) begin
      lineBuffer_321 <= lineBuffer_320;
    end
    if (sel) begin
      lineBuffer_322 <= lineBuffer_321;
    end
    if (sel) begin
      lineBuffer_323 <= lineBuffer_322;
    end
    if (sel) begin
      lineBuffer_324 <= lineBuffer_323;
    end
    if (sel) begin
      lineBuffer_325 <= lineBuffer_324;
    end
    if (sel) begin
      lineBuffer_326 <= lineBuffer_325;
    end
    if (sel) begin
      lineBuffer_327 <= lineBuffer_326;
    end
    if (sel) begin
      lineBuffer_328 <= lineBuffer_327;
    end
    if (sel) begin
      lineBuffer_329 <= lineBuffer_328;
    end
    if (sel) begin
      lineBuffer_330 <= lineBuffer_329;
    end
    if (sel) begin
      lineBuffer_331 <= lineBuffer_330;
    end
    if (sel) begin
      lineBuffer_332 <= lineBuffer_331;
    end
    if (sel) begin
      lineBuffer_333 <= lineBuffer_332;
    end
    if (sel) begin
      lineBuffer_334 <= lineBuffer_333;
    end
    if (sel) begin
      lineBuffer_335 <= lineBuffer_334;
    end
    if (sel) begin
      lineBuffer_336 <= lineBuffer_335;
    end
    if (sel) begin
      lineBuffer_337 <= lineBuffer_336;
    end
    if (sel) begin
      lineBuffer_338 <= lineBuffer_337;
    end
    if (sel) begin
      lineBuffer_339 <= lineBuffer_338;
    end
    if (sel) begin
      lineBuffer_340 <= lineBuffer_339;
    end
    if (sel) begin
      lineBuffer_341 <= lineBuffer_340;
    end
    if (sel) begin
      lineBuffer_342 <= lineBuffer_341;
    end
    if (sel) begin
      lineBuffer_343 <= lineBuffer_342;
    end
    if (sel) begin
      lineBuffer_344 <= lineBuffer_343;
    end
    if (sel) begin
      lineBuffer_345 <= lineBuffer_344;
    end
    if (sel) begin
      lineBuffer_346 <= lineBuffer_345;
    end
    if (sel) begin
      lineBuffer_347 <= lineBuffer_346;
    end
    if (sel) begin
      lineBuffer_348 <= lineBuffer_347;
    end
    if (sel) begin
      lineBuffer_349 <= lineBuffer_348;
    end
    if (sel) begin
      lineBuffer_350 <= lineBuffer_349;
    end
    if (sel) begin
      lineBuffer_351 <= lineBuffer_350;
    end
    if (sel) begin
      lineBuffer_352 <= lineBuffer_351;
    end
    if (sel) begin
      lineBuffer_353 <= lineBuffer_352;
    end
    if (sel) begin
      lineBuffer_354 <= lineBuffer_353;
    end
    if (sel) begin
      lineBuffer_355 <= lineBuffer_354;
    end
    if (sel) begin
      lineBuffer_356 <= lineBuffer_355;
    end
    if (sel) begin
      lineBuffer_357 <= lineBuffer_356;
    end
    if (sel) begin
      lineBuffer_358 <= lineBuffer_357;
    end
    if (sel) begin
      lineBuffer_359 <= lineBuffer_358;
    end
    if (sel) begin
      lineBuffer_360 <= lineBuffer_359;
    end
    if (sel) begin
      lineBuffer_361 <= lineBuffer_360;
    end
    if (sel) begin
      lineBuffer_362 <= lineBuffer_361;
    end
    if (sel) begin
      lineBuffer_363 <= lineBuffer_362;
    end
    if (sel) begin
      lineBuffer_364 <= lineBuffer_363;
    end
    if (sel) begin
      lineBuffer_365 <= lineBuffer_364;
    end
    if (sel) begin
      lineBuffer_366 <= lineBuffer_365;
    end
    if (sel) begin
      lineBuffer_367 <= lineBuffer_366;
    end
    if (sel) begin
      lineBuffer_368 <= lineBuffer_367;
    end
    if (sel) begin
      lineBuffer_369 <= lineBuffer_368;
    end
    if (sel) begin
      lineBuffer_370 <= lineBuffer_369;
    end
    if (sel) begin
      lineBuffer_371 <= lineBuffer_370;
    end
    if (sel) begin
      lineBuffer_372 <= lineBuffer_371;
    end
    if (sel) begin
      lineBuffer_373 <= lineBuffer_372;
    end
    if (sel) begin
      lineBuffer_374 <= lineBuffer_373;
    end
    if (sel) begin
      lineBuffer_375 <= lineBuffer_374;
    end
    if (sel) begin
      lineBuffer_376 <= lineBuffer_375;
    end
    if (sel) begin
      lineBuffer_377 <= lineBuffer_376;
    end
    if (sel) begin
      lineBuffer_378 <= lineBuffer_377;
    end
    if (sel) begin
      lineBuffer_379 <= lineBuffer_378;
    end
    if (sel) begin
      lineBuffer_380 <= lineBuffer_379;
    end
    if (sel) begin
      lineBuffer_381 <= lineBuffer_380;
    end
    if (sel) begin
      lineBuffer_382 <= lineBuffer_381;
    end
    if (sel) begin
      lineBuffer_383 <= lineBuffer_382;
    end
    if (sel) begin
      lineBuffer_384 <= lineBuffer_383;
    end
    if (sel) begin
      lineBuffer_385 <= lineBuffer_384;
    end
    if (sel) begin
      lineBuffer_386 <= lineBuffer_385;
    end
    if (sel) begin
      lineBuffer_387 <= lineBuffer_386;
    end
    if (sel) begin
      lineBuffer_388 <= lineBuffer_387;
    end
    if (sel) begin
      lineBuffer_389 <= lineBuffer_388;
    end
    if (sel) begin
      lineBuffer_390 <= lineBuffer_389;
    end
    if (sel) begin
      lineBuffer_391 <= lineBuffer_390;
    end
    if (sel) begin
      lineBuffer_392 <= lineBuffer_391;
    end
    if (sel) begin
      lineBuffer_393 <= lineBuffer_392;
    end
    if (sel) begin
      lineBuffer_394 <= lineBuffer_393;
    end
    if (sel) begin
      lineBuffer_395 <= lineBuffer_394;
    end
    if (sel) begin
      lineBuffer_396 <= lineBuffer_395;
    end
    if (sel) begin
      lineBuffer_397 <= lineBuffer_396;
    end
    if (sel) begin
      lineBuffer_398 <= lineBuffer_397;
    end
    if (sel) begin
      lineBuffer_399 <= lineBuffer_398;
    end
    if (sel) begin
      lineBuffer_400 <= lineBuffer_399;
    end
    if (sel) begin
      lineBuffer_401 <= lineBuffer_400;
    end
    if (sel) begin
      lineBuffer_402 <= lineBuffer_401;
    end
    if (sel) begin
      lineBuffer_403 <= lineBuffer_402;
    end
    if (sel) begin
      lineBuffer_404 <= lineBuffer_403;
    end
    if (sel) begin
      lineBuffer_405 <= lineBuffer_404;
    end
    if (sel) begin
      lineBuffer_406 <= lineBuffer_405;
    end
    if (sel) begin
      lineBuffer_407 <= lineBuffer_406;
    end
    if (sel) begin
      lineBuffer_408 <= lineBuffer_407;
    end
    if (sel) begin
      lineBuffer_409 <= lineBuffer_408;
    end
    if (sel) begin
      lineBuffer_410 <= lineBuffer_409;
    end
    if (sel) begin
      lineBuffer_411 <= lineBuffer_410;
    end
    if (sel) begin
      lineBuffer_412 <= lineBuffer_411;
    end
    if (sel) begin
      lineBuffer_413 <= lineBuffer_412;
    end
    if (sel) begin
      lineBuffer_414 <= lineBuffer_413;
    end
    if (sel) begin
      lineBuffer_415 <= lineBuffer_414;
    end
    if (sel) begin
      lineBuffer_416 <= lineBuffer_415;
    end
    if (sel) begin
      lineBuffer_417 <= lineBuffer_416;
    end
    if (sel) begin
      lineBuffer_418 <= lineBuffer_417;
    end
    if (sel) begin
      lineBuffer_419 <= lineBuffer_418;
    end
    if (sel) begin
      lineBuffer_420 <= lineBuffer_419;
    end
    if (sel) begin
      lineBuffer_421 <= lineBuffer_420;
    end
    if (sel) begin
      lineBuffer_422 <= lineBuffer_421;
    end
    if (sel) begin
      lineBuffer_423 <= lineBuffer_422;
    end
    if (sel) begin
      lineBuffer_424 <= lineBuffer_423;
    end
    if (sel) begin
      lineBuffer_425 <= lineBuffer_424;
    end
    if (sel) begin
      lineBuffer_426 <= lineBuffer_425;
    end
    if (sel) begin
      lineBuffer_427 <= lineBuffer_426;
    end
    if (sel) begin
      lineBuffer_428 <= lineBuffer_427;
    end
    if (sel) begin
      lineBuffer_429 <= lineBuffer_428;
    end
    if (sel) begin
      lineBuffer_430 <= lineBuffer_429;
    end
    if (sel) begin
      lineBuffer_431 <= lineBuffer_430;
    end
    if (sel) begin
      lineBuffer_432 <= lineBuffer_431;
    end
    if (sel) begin
      lineBuffer_433 <= lineBuffer_432;
    end
    if (sel) begin
      lineBuffer_434 <= lineBuffer_433;
    end
    if (sel) begin
      lineBuffer_435 <= lineBuffer_434;
    end
    if (sel) begin
      lineBuffer_436 <= lineBuffer_435;
    end
    if (sel) begin
      lineBuffer_437 <= lineBuffer_436;
    end
    if (sel) begin
      lineBuffer_438 <= lineBuffer_437;
    end
    if (sel) begin
      lineBuffer_439 <= lineBuffer_438;
    end
    if (sel) begin
      lineBuffer_440 <= lineBuffer_439;
    end
    if (sel) begin
      lineBuffer_441 <= lineBuffer_440;
    end
    if (sel) begin
      lineBuffer_442 <= lineBuffer_441;
    end
    if (sel) begin
      lineBuffer_443 <= lineBuffer_442;
    end
    if (sel) begin
      lineBuffer_444 <= lineBuffer_443;
    end
    if (sel) begin
      lineBuffer_445 <= lineBuffer_444;
    end
    if (sel) begin
      lineBuffer_446 <= lineBuffer_445;
    end
    if (sel) begin
      lineBuffer_447 <= lineBuffer_446;
    end
    if (sel) begin
      lineBuffer_448 <= lineBuffer_447;
    end
    if (sel) begin
      lineBuffer_449 <= lineBuffer_448;
    end
    if (sel) begin
      lineBuffer_450 <= lineBuffer_449;
    end
    if (sel) begin
      lineBuffer_451 <= lineBuffer_450;
    end
    if (sel) begin
      lineBuffer_452 <= lineBuffer_451;
    end
    if (sel) begin
      lineBuffer_453 <= lineBuffer_452;
    end
    if (sel) begin
      lineBuffer_454 <= lineBuffer_453;
    end
    if (sel) begin
      lineBuffer_455 <= lineBuffer_454;
    end
    if (sel) begin
      lineBuffer_456 <= lineBuffer_455;
    end
    if (sel) begin
      lineBuffer_457 <= lineBuffer_456;
    end
    if (sel) begin
      lineBuffer_458 <= lineBuffer_457;
    end
    if (sel) begin
      lineBuffer_459 <= lineBuffer_458;
    end
    if (sel) begin
      lineBuffer_460 <= lineBuffer_459;
    end
    if (sel) begin
      lineBuffer_461 <= lineBuffer_460;
    end
    if (sel) begin
      lineBuffer_462 <= lineBuffer_461;
    end
    if (sel) begin
      lineBuffer_463 <= lineBuffer_462;
    end
    if (sel) begin
      lineBuffer_464 <= lineBuffer_463;
    end
    if (sel) begin
      lineBuffer_465 <= lineBuffer_464;
    end
    if (sel) begin
      lineBuffer_466 <= lineBuffer_465;
    end
    if (sel) begin
      lineBuffer_467 <= lineBuffer_466;
    end
    if (sel) begin
      lineBuffer_468 <= lineBuffer_467;
    end
    if (sel) begin
      lineBuffer_469 <= lineBuffer_468;
    end
    if (sel) begin
      lineBuffer_470 <= lineBuffer_469;
    end
    if (sel) begin
      lineBuffer_471 <= lineBuffer_470;
    end
    if (sel) begin
      lineBuffer_472 <= lineBuffer_471;
    end
    if (sel) begin
      lineBuffer_473 <= lineBuffer_472;
    end
    if (sel) begin
      lineBuffer_474 <= lineBuffer_473;
    end
    if (sel) begin
      lineBuffer_475 <= lineBuffer_474;
    end
    if (sel) begin
      lineBuffer_476 <= lineBuffer_475;
    end
    if (sel) begin
      lineBuffer_477 <= lineBuffer_476;
    end
    if (sel) begin
      lineBuffer_478 <= lineBuffer_477;
    end
    if (sel) begin
      lineBuffer_479 <= lineBuffer_478;
    end
    if (sel) begin
      lineBuffer_480 <= lineBuffer_479;
    end
    if (sel) begin
      lineBuffer_481 <= lineBuffer_480;
    end
    if (sel) begin
      lineBuffer_482 <= lineBuffer_481;
    end
    if (sel) begin
      lineBuffer_483 <= lineBuffer_482;
    end
    if (sel) begin
      lineBuffer_484 <= lineBuffer_483;
    end
    if (sel) begin
      lineBuffer_485 <= lineBuffer_484;
    end
    if (sel) begin
      lineBuffer_486 <= lineBuffer_485;
    end
    if (sel) begin
      lineBuffer_487 <= lineBuffer_486;
    end
    if (sel) begin
      lineBuffer_488 <= lineBuffer_487;
    end
    if (sel) begin
      lineBuffer_489 <= lineBuffer_488;
    end
    if (sel) begin
      lineBuffer_490 <= lineBuffer_489;
    end
    if (sel) begin
      lineBuffer_491 <= lineBuffer_490;
    end
    if (sel) begin
      lineBuffer_492 <= lineBuffer_491;
    end
    if (sel) begin
      lineBuffer_493 <= lineBuffer_492;
    end
    if (sel) begin
      lineBuffer_494 <= lineBuffer_493;
    end
    if (sel) begin
      lineBuffer_495 <= lineBuffer_494;
    end
    if (sel) begin
      lineBuffer_496 <= lineBuffer_495;
    end
    if (sel) begin
      lineBuffer_497 <= lineBuffer_496;
    end
    if (sel) begin
      lineBuffer_498 <= lineBuffer_497;
    end
    if (sel) begin
      lineBuffer_499 <= lineBuffer_498;
    end
    if (sel) begin
      lineBuffer_500 <= lineBuffer_499;
    end
    if (sel) begin
      lineBuffer_501 <= lineBuffer_500;
    end
    if (sel) begin
      lineBuffer_502 <= lineBuffer_501;
    end
    if (sel) begin
      lineBuffer_503 <= lineBuffer_502;
    end
    if (sel) begin
      lineBuffer_504 <= lineBuffer_503;
    end
    if (sel) begin
      lineBuffer_505 <= lineBuffer_504;
    end
    if (sel) begin
      lineBuffer_506 <= lineBuffer_505;
    end
    if (sel) begin
      lineBuffer_507 <= lineBuffer_506;
    end
    if (sel) begin
      lineBuffer_508 <= lineBuffer_507;
    end
    if (sel) begin
      lineBuffer_509 <= lineBuffer_508;
    end
    if (sel) begin
      lineBuffer_510 <= lineBuffer_509;
    end
    if (sel) begin
      lineBuffer_511 <= lineBuffer_510;
    end
    if (sel) begin
      lineBuffer_512 <= lineBuffer_511;
    end
    if (sel) begin
      lineBuffer_513 <= lineBuffer_512;
    end
    if (sel) begin
      lineBuffer_514 <= lineBuffer_513;
    end
    if (sel) begin
      lineBuffer_515 <= lineBuffer_514;
    end
    if (sel) begin
      lineBuffer_516 <= lineBuffer_515;
    end
    if (sel) begin
      lineBuffer_517 <= lineBuffer_516;
    end
    if (sel) begin
      lineBuffer_518 <= lineBuffer_517;
    end
    if (sel) begin
      lineBuffer_519 <= lineBuffer_518;
    end
    if (sel) begin
      lineBuffer_520 <= lineBuffer_519;
    end
    if (sel) begin
      lineBuffer_521 <= lineBuffer_520;
    end
    if (sel) begin
      lineBuffer_522 <= lineBuffer_521;
    end
    if (sel) begin
      lineBuffer_523 <= lineBuffer_522;
    end
    if (sel) begin
      lineBuffer_524 <= lineBuffer_523;
    end
    if (sel) begin
      lineBuffer_525 <= lineBuffer_524;
    end
    if (sel) begin
      lineBuffer_526 <= lineBuffer_525;
    end
    if (sel) begin
      lineBuffer_527 <= lineBuffer_526;
    end
    if (sel) begin
      lineBuffer_528 <= lineBuffer_527;
    end
    if (sel) begin
      lineBuffer_529 <= lineBuffer_528;
    end
    if (sel) begin
      lineBuffer_530 <= lineBuffer_529;
    end
    if (sel) begin
      lineBuffer_531 <= lineBuffer_530;
    end
    if (sel) begin
      lineBuffer_532 <= lineBuffer_531;
    end
    if (sel) begin
      lineBuffer_533 <= lineBuffer_532;
    end
    if (sel) begin
      lineBuffer_534 <= lineBuffer_533;
    end
    if (sel) begin
      lineBuffer_535 <= lineBuffer_534;
    end
    if (sel) begin
      lineBuffer_536 <= lineBuffer_535;
    end
    if (sel) begin
      lineBuffer_537 <= lineBuffer_536;
    end
    if (sel) begin
      lineBuffer_538 <= lineBuffer_537;
    end
    if (sel) begin
      lineBuffer_539 <= lineBuffer_538;
    end
    if (sel) begin
      lineBuffer_540 <= lineBuffer_539;
    end
    if (sel) begin
      lineBuffer_541 <= lineBuffer_540;
    end
    if (sel) begin
      lineBuffer_542 <= lineBuffer_541;
    end
    if (sel) begin
      lineBuffer_543 <= lineBuffer_542;
    end
    if (sel) begin
      lineBuffer_544 <= lineBuffer_543;
    end
    if (sel) begin
      lineBuffer_545 <= lineBuffer_544;
    end
    if (sel) begin
      lineBuffer_546 <= lineBuffer_545;
    end
    if (sel) begin
      lineBuffer_547 <= lineBuffer_546;
    end
    if (sel) begin
      lineBuffer_548 <= lineBuffer_547;
    end
    if (sel) begin
      lineBuffer_549 <= lineBuffer_548;
    end
    if (sel) begin
      lineBuffer_550 <= lineBuffer_549;
    end
    if (sel) begin
      lineBuffer_551 <= lineBuffer_550;
    end
    if (sel) begin
      lineBuffer_552 <= lineBuffer_551;
    end
    if (sel) begin
      lineBuffer_553 <= lineBuffer_552;
    end
    if (sel) begin
      lineBuffer_554 <= lineBuffer_553;
    end
    if (sel) begin
      lineBuffer_555 <= lineBuffer_554;
    end
    if (sel) begin
      lineBuffer_556 <= lineBuffer_555;
    end
    if (sel) begin
      lineBuffer_557 <= lineBuffer_556;
    end
    if (sel) begin
      lineBuffer_558 <= lineBuffer_557;
    end
    if (sel) begin
      lineBuffer_559 <= lineBuffer_558;
    end
    if (sel) begin
      lineBuffer_560 <= lineBuffer_559;
    end
    if (sel) begin
      lineBuffer_561 <= lineBuffer_560;
    end
    if (sel) begin
      lineBuffer_562 <= lineBuffer_561;
    end
    if (sel) begin
      lineBuffer_563 <= lineBuffer_562;
    end
    if (sel) begin
      lineBuffer_564 <= lineBuffer_563;
    end
    if (sel) begin
      lineBuffer_565 <= lineBuffer_564;
    end
    if (sel) begin
      lineBuffer_566 <= lineBuffer_565;
    end
    if (sel) begin
      lineBuffer_567 <= lineBuffer_566;
    end
    if (sel) begin
      lineBuffer_568 <= lineBuffer_567;
    end
    if (sel) begin
      lineBuffer_569 <= lineBuffer_568;
    end
    if (sel) begin
      lineBuffer_570 <= lineBuffer_569;
    end
    if (sel) begin
      lineBuffer_571 <= lineBuffer_570;
    end
    if (sel) begin
      lineBuffer_572 <= lineBuffer_571;
    end
    if (sel) begin
      lineBuffer_573 <= lineBuffer_572;
    end
    if (sel) begin
      lineBuffer_574 <= lineBuffer_573;
    end
    if (sel) begin
      lineBuffer_575 <= lineBuffer_574;
    end
    if (sel) begin
      lineBuffer_576 <= lineBuffer_575;
    end
    if (sel) begin
      lineBuffer_577 <= lineBuffer_576;
    end
    if (sel) begin
      lineBuffer_578 <= lineBuffer_577;
    end
    if (sel) begin
      lineBuffer_579 <= lineBuffer_578;
    end
    if (sel) begin
      lineBuffer_580 <= lineBuffer_579;
    end
    if (sel) begin
      lineBuffer_581 <= lineBuffer_580;
    end
    if (sel) begin
      lineBuffer_582 <= lineBuffer_581;
    end
    if (sel) begin
      lineBuffer_583 <= lineBuffer_582;
    end
    if (sel) begin
      lineBuffer_584 <= lineBuffer_583;
    end
    if (sel) begin
      lineBuffer_585 <= lineBuffer_584;
    end
    if (sel) begin
      lineBuffer_586 <= lineBuffer_585;
    end
    if (sel) begin
      lineBuffer_587 <= lineBuffer_586;
    end
    if (sel) begin
      lineBuffer_588 <= lineBuffer_587;
    end
    if (sel) begin
      lineBuffer_589 <= lineBuffer_588;
    end
    if (sel) begin
      lineBuffer_590 <= lineBuffer_589;
    end
    if (sel) begin
      lineBuffer_591 <= lineBuffer_590;
    end
    if (sel) begin
      lineBuffer_592 <= lineBuffer_591;
    end
    if (sel) begin
      lineBuffer_593 <= lineBuffer_592;
    end
    if (sel) begin
      lineBuffer_594 <= lineBuffer_593;
    end
    if (sel) begin
      lineBuffer_595 <= lineBuffer_594;
    end
    if (sel) begin
      lineBuffer_596 <= lineBuffer_595;
    end
    if (sel) begin
      lineBuffer_597 <= lineBuffer_596;
    end
    if (sel) begin
      lineBuffer_598 <= lineBuffer_597;
    end
    if (sel) begin
      lineBuffer_599 <= lineBuffer_598;
    end
    if (sel) begin
      lineBuffer_600 <= lineBuffer_599;
    end
    if (sel) begin
      lineBuffer_601 <= lineBuffer_600;
    end
    if (sel) begin
      lineBuffer_602 <= lineBuffer_601;
    end
    if (sel) begin
      lineBuffer_603 <= lineBuffer_602;
    end
    if (sel) begin
      lineBuffer_604 <= lineBuffer_603;
    end
    if (sel) begin
      lineBuffer_605 <= lineBuffer_604;
    end
    if (sel) begin
      lineBuffer_606 <= lineBuffer_605;
    end
    if (sel) begin
      lineBuffer_607 <= lineBuffer_606;
    end
    if (sel) begin
      lineBuffer_608 <= lineBuffer_607;
    end
    if (sel) begin
      lineBuffer_609 <= lineBuffer_608;
    end
    if (sel) begin
      lineBuffer_610 <= lineBuffer_609;
    end
    if (sel) begin
      lineBuffer_611 <= lineBuffer_610;
    end
    if (sel) begin
      lineBuffer_612 <= lineBuffer_611;
    end
    if (sel) begin
      lineBuffer_613 <= lineBuffer_612;
    end
    if (sel) begin
      lineBuffer_614 <= lineBuffer_613;
    end
    if (sel) begin
      lineBuffer_615 <= lineBuffer_614;
    end
    if (sel) begin
      lineBuffer_616 <= lineBuffer_615;
    end
    if (sel) begin
      lineBuffer_617 <= lineBuffer_616;
    end
    if (sel) begin
      lineBuffer_618 <= lineBuffer_617;
    end
    if (sel) begin
      lineBuffer_619 <= lineBuffer_618;
    end
    if (sel) begin
      lineBuffer_620 <= lineBuffer_619;
    end
    if (sel) begin
      lineBuffer_621 <= lineBuffer_620;
    end
    if (sel) begin
      lineBuffer_622 <= lineBuffer_621;
    end
    if (sel) begin
      lineBuffer_623 <= lineBuffer_622;
    end
    if (sel) begin
      lineBuffer_624 <= lineBuffer_623;
    end
    if (sel) begin
      lineBuffer_625 <= lineBuffer_624;
    end
    if (sel) begin
      lineBuffer_626 <= lineBuffer_625;
    end
    if (sel) begin
      lineBuffer_627 <= lineBuffer_626;
    end
    if (sel) begin
      lineBuffer_628 <= lineBuffer_627;
    end
    if (sel) begin
      lineBuffer_629 <= lineBuffer_628;
    end
    if (sel) begin
      lineBuffer_630 <= lineBuffer_629;
    end
    if (sel) begin
      lineBuffer_631 <= lineBuffer_630;
    end
    if (sel) begin
      lineBuffer_632 <= lineBuffer_631;
    end
    if (sel) begin
      lineBuffer_633 <= lineBuffer_632;
    end
    if (sel) begin
      lineBuffer_634 <= lineBuffer_633;
    end
    if (sel) begin
      lineBuffer_635 <= lineBuffer_634;
    end
    if (sel) begin
      lineBuffer_636 <= lineBuffer_635;
    end
    if (sel) begin
      lineBuffer_637 <= lineBuffer_636;
    end
    if (sel) begin
      lineBuffer_638 <= lineBuffer_637;
    end
    if (sel) begin
      lineBuffer_639 <= lineBuffer_638;
    end
    if (sel) begin
      lineBuffer_640 <= lineBuffer_639;
    end
    if (sel) begin
      lineBuffer_641 <= lineBuffer_640;
    end
    if (sel) begin
      lineBuffer_642 <= lineBuffer_641;
    end
    if (sel) begin
      lineBuffer_643 <= lineBuffer_642;
    end
    if (sel) begin
      lineBuffer_644 <= lineBuffer_643;
    end
    if (sel) begin
      lineBuffer_645 <= lineBuffer_644;
    end
    if (sel) begin
      lineBuffer_646 <= lineBuffer_645;
    end
    if (sel) begin
      lineBuffer_647 <= lineBuffer_646;
    end
    if (sel) begin
      lineBuffer_648 <= lineBuffer_647;
    end
    if (sel) begin
      lineBuffer_649 <= lineBuffer_648;
    end
    if (sel) begin
      lineBuffer_650 <= lineBuffer_649;
    end
    if (sel) begin
      lineBuffer_651 <= lineBuffer_650;
    end
    if (sel) begin
      lineBuffer_652 <= lineBuffer_651;
    end
    if (sel) begin
      lineBuffer_653 <= lineBuffer_652;
    end
    if (sel) begin
      lineBuffer_654 <= lineBuffer_653;
    end
    if (sel) begin
      lineBuffer_655 <= lineBuffer_654;
    end
    if (sel) begin
      lineBuffer_656 <= lineBuffer_655;
    end
    if (sel) begin
      lineBuffer_657 <= lineBuffer_656;
    end
    if (sel) begin
      lineBuffer_658 <= lineBuffer_657;
    end
    if (sel) begin
      lineBuffer_659 <= lineBuffer_658;
    end
    if (sel) begin
      lineBuffer_660 <= lineBuffer_659;
    end
    if (sel) begin
      lineBuffer_661 <= lineBuffer_660;
    end
    if (sel) begin
      lineBuffer_662 <= lineBuffer_661;
    end
    if (sel) begin
      lineBuffer_663 <= lineBuffer_662;
    end
    if (sel) begin
      lineBuffer_664 <= lineBuffer_663;
    end
    if (sel) begin
      lineBuffer_665 <= lineBuffer_664;
    end
    if (sel) begin
      lineBuffer_666 <= lineBuffer_665;
    end
    if (sel) begin
      lineBuffer_667 <= lineBuffer_666;
    end
    if (sel) begin
      lineBuffer_668 <= lineBuffer_667;
    end
    if (sel) begin
      lineBuffer_669 <= lineBuffer_668;
    end
    if (sel) begin
      lineBuffer_670 <= lineBuffer_669;
    end
    if (sel) begin
      lineBuffer_671 <= lineBuffer_670;
    end
    if (sel) begin
      lineBuffer_672 <= lineBuffer_671;
    end
    if (sel) begin
      lineBuffer_673 <= lineBuffer_672;
    end
    if (sel) begin
      lineBuffer_674 <= lineBuffer_673;
    end
    if (sel) begin
      lineBuffer_675 <= lineBuffer_674;
    end
    if (sel) begin
      lineBuffer_676 <= lineBuffer_675;
    end
    if (sel) begin
      lineBuffer_677 <= lineBuffer_676;
    end
    if (sel) begin
      lineBuffer_678 <= lineBuffer_677;
    end
    if (sel) begin
      lineBuffer_679 <= lineBuffer_678;
    end
    if (sel) begin
      lineBuffer_680 <= lineBuffer_679;
    end
    if (sel) begin
      lineBuffer_681 <= lineBuffer_680;
    end
    if (sel) begin
      lineBuffer_682 <= lineBuffer_681;
    end
    if (sel) begin
      lineBuffer_683 <= lineBuffer_682;
    end
    if (sel) begin
      lineBuffer_684 <= lineBuffer_683;
    end
    if (sel) begin
      lineBuffer_685 <= lineBuffer_684;
    end
    if (sel) begin
      lineBuffer_686 <= lineBuffer_685;
    end
    if (sel) begin
      lineBuffer_687 <= lineBuffer_686;
    end
    if (sel) begin
      lineBuffer_688 <= lineBuffer_687;
    end
    if (sel) begin
      lineBuffer_689 <= lineBuffer_688;
    end
    if (sel) begin
      lineBuffer_690 <= lineBuffer_689;
    end
    if (sel) begin
      lineBuffer_691 <= lineBuffer_690;
    end
    if (sel) begin
      lineBuffer_692 <= lineBuffer_691;
    end
    if (sel) begin
      lineBuffer_693 <= lineBuffer_692;
    end
    if (sel) begin
      lineBuffer_694 <= lineBuffer_693;
    end
    if (sel) begin
      lineBuffer_695 <= lineBuffer_694;
    end
    if (sel) begin
      lineBuffer_696 <= lineBuffer_695;
    end
    if (sel) begin
      lineBuffer_697 <= lineBuffer_696;
    end
    if (sel) begin
      lineBuffer_698 <= lineBuffer_697;
    end
    if (sel) begin
      lineBuffer_699 <= lineBuffer_698;
    end
    if (sel) begin
      lineBuffer_700 <= lineBuffer_699;
    end
    if (sel) begin
      lineBuffer_701 <= lineBuffer_700;
    end
    if (sel) begin
      lineBuffer_702 <= lineBuffer_701;
    end
    if (sel) begin
      lineBuffer_703 <= lineBuffer_702;
    end
    if (sel) begin
      lineBuffer_704 <= lineBuffer_703;
    end
    if (sel) begin
      lineBuffer_705 <= lineBuffer_704;
    end
    if (sel) begin
      lineBuffer_706 <= lineBuffer_705;
    end
    if (sel) begin
      lineBuffer_707 <= lineBuffer_706;
    end
    if (sel) begin
      lineBuffer_708 <= lineBuffer_707;
    end
    if (sel) begin
      lineBuffer_709 <= lineBuffer_708;
    end
    if (sel) begin
      lineBuffer_710 <= lineBuffer_709;
    end
    if (sel) begin
      lineBuffer_711 <= lineBuffer_710;
    end
    if (sel) begin
      lineBuffer_712 <= lineBuffer_711;
    end
    if (sel) begin
      lineBuffer_713 <= lineBuffer_712;
    end
    if (sel) begin
      lineBuffer_714 <= lineBuffer_713;
    end
    if (sel) begin
      lineBuffer_715 <= lineBuffer_714;
    end
    if (sel) begin
      lineBuffer_716 <= lineBuffer_715;
    end
    if (sel) begin
      lineBuffer_717 <= lineBuffer_716;
    end
    if (sel) begin
      lineBuffer_718 <= lineBuffer_717;
    end
    if (sel) begin
      lineBuffer_719 <= lineBuffer_718;
    end
    if (sel) begin
      lineBuffer_720 <= lineBuffer_719;
    end
    if (sel) begin
      lineBuffer_721 <= lineBuffer_720;
    end
    if (sel) begin
      lineBuffer_722 <= lineBuffer_721;
    end
    if (sel) begin
      lineBuffer_723 <= lineBuffer_722;
    end
    if (sel) begin
      lineBuffer_724 <= lineBuffer_723;
    end
    if (sel) begin
      lineBuffer_725 <= lineBuffer_724;
    end
    if (sel) begin
      lineBuffer_726 <= lineBuffer_725;
    end
    if (sel) begin
      lineBuffer_727 <= lineBuffer_726;
    end
    if (sel) begin
      lineBuffer_728 <= lineBuffer_727;
    end
    if (sel) begin
      lineBuffer_729 <= lineBuffer_728;
    end
    if (sel) begin
      lineBuffer_730 <= lineBuffer_729;
    end
    if (sel) begin
      lineBuffer_731 <= lineBuffer_730;
    end
    if (sel) begin
      lineBuffer_732 <= lineBuffer_731;
    end
    if (sel) begin
      lineBuffer_733 <= lineBuffer_732;
    end
    if (sel) begin
      lineBuffer_734 <= lineBuffer_733;
    end
    if (sel) begin
      lineBuffer_735 <= lineBuffer_734;
    end
    if (sel) begin
      lineBuffer_736 <= lineBuffer_735;
    end
    if (sel) begin
      lineBuffer_737 <= lineBuffer_736;
    end
    if (sel) begin
      lineBuffer_738 <= lineBuffer_737;
    end
    if (sel) begin
      lineBuffer_739 <= lineBuffer_738;
    end
    if (sel) begin
      lineBuffer_740 <= lineBuffer_739;
    end
    if (sel) begin
      lineBuffer_741 <= lineBuffer_740;
    end
    if (sel) begin
      lineBuffer_742 <= lineBuffer_741;
    end
    if (sel) begin
      lineBuffer_743 <= lineBuffer_742;
    end
    if (sel) begin
      lineBuffer_744 <= lineBuffer_743;
    end
    if (sel) begin
      lineBuffer_745 <= lineBuffer_744;
    end
    if (sel) begin
      lineBuffer_746 <= lineBuffer_745;
    end
    if (sel) begin
      lineBuffer_747 <= lineBuffer_746;
    end
    if (sel) begin
      lineBuffer_748 <= lineBuffer_747;
    end
    if (sel) begin
      lineBuffer_749 <= lineBuffer_748;
    end
    if (sel) begin
      lineBuffer_750 <= lineBuffer_749;
    end
    if (sel) begin
      lineBuffer_751 <= lineBuffer_750;
    end
    if (sel) begin
      lineBuffer_752 <= lineBuffer_751;
    end
    if (sel) begin
      lineBuffer_753 <= lineBuffer_752;
    end
    if (sel) begin
      lineBuffer_754 <= lineBuffer_753;
    end
    if (sel) begin
      lineBuffer_755 <= lineBuffer_754;
    end
    if (sel) begin
      lineBuffer_756 <= lineBuffer_755;
    end
    if (sel) begin
      lineBuffer_757 <= lineBuffer_756;
    end
    if (sel) begin
      lineBuffer_758 <= lineBuffer_757;
    end
    if (sel) begin
      lineBuffer_759 <= lineBuffer_758;
    end
    if (sel) begin
      lineBuffer_760 <= lineBuffer_759;
    end
    if (sel) begin
      lineBuffer_761 <= lineBuffer_760;
    end
    if (sel) begin
      lineBuffer_762 <= lineBuffer_761;
    end
    if (sel) begin
      lineBuffer_763 <= lineBuffer_762;
    end
    if (sel) begin
      lineBuffer_764 <= lineBuffer_763;
    end
    if (sel) begin
      lineBuffer_765 <= lineBuffer_764;
    end
    if (sel) begin
      lineBuffer_766 <= lineBuffer_765;
    end
    if (sel) begin
      lineBuffer_767 <= lineBuffer_766;
    end
    if (sel) begin
      windowBuffer_0 <= windowBuffer_1;
    end
    if (sel) begin
      windowBuffer_1 <= windowBuffer_2;
    end
    if (sel) begin
      windowBuffer_2 <= lineBuffer_255;
    end
    if (sel) begin
      windowBuffer_3 <= windowBuffer_4;
    end
    if (sel) begin
      windowBuffer_4 <= windowBuffer_5;
    end
    if (sel) begin
      windowBuffer_5 <= lineBuffer_511;
    end
    if (sel) begin
      windowBuffer_6 <= windowBuffer_7;
    end
    if (sel) begin
      windowBuffer_7 <= windowBuffer_8;
    end
    if (sel) begin
      windowBuffer_8 <= lineBuffer_767;
    end
  end
endmodule
module SMulAdd(
  input  [15:0] io_a_1,
  input  [15:0] io_a_2,
  input  [15:0] io_a_3,
  input  [15:0] io_a_5,
  input  [15:0] io_a_6,
  input  [15:0] io_a_7,
  input  [15:0] io_b_0,
  input  [15:0] io_b_1,
  input  [15:0] io_b_2,
  input  [15:0] io_b_3,
  input  [15:0] io_b_4,
  input  [15:0] io_b_5,
  input  [15:0] io_b_6,
  input  [15:0] io_b_7,
  input  [15:0] io_b_8,
  output [31:0] io_output
);
  wire [31:0] _T = 16'sh1 * $signed(io_b_0); // @[ChiselImProc.scala 50:24]
  wire [32:0] _T_1 = {{1{_T[31]}},_T}; // @[ChiselImProc.scala 50:13]
  wire [31:0] _T_3 = _T_1[31:0]; // @[ChiselImProc.scala 50:13]
  wire [31:0] _T_4 = $signed(io_a_1) * $signed(io_b_1); // @[ChiselImProc.scala 50:24]
  wire [31:0] _T_7 = $signed(_T_3) + $signed(_T_4); // @[ChiselImProc.scala 50:13]
  wire [31:0] _T_8 = $signed(io_a_2) * $signed(io_b_2); // @[ChiselImProc.scala 50:24]
  wire [31:0] _T_11 = $signed(_T_7) + $signed(_T_8); // @[ChiselImProc.scala 50:13]
  wire [31:0] _T_12 = $signed(io_a_3) * $signed(io_b_3); // @[ChiselImProc.scala 50:24]
  wire [31:0] _T_15 = $signed(_T_11) + $signed(_T_12); // @[ChiselImProc.scala 50:13]
  wire [31:0] _T_16 = 16'sh0 * $signed(io_b_4); // @[ChiselImProc.scala 50:24]
  wire [31:0] _T_19 = $signed(_T_15) + $signed(_T_16); // @[ChiselImProc.scala 50:13]
  wire [31:0] _T_20 = $signed(io_a_5) * $signed(io_b_5); // @[ChiselImProc.scala 50:24]
  wire [31:0] _T_23 = $signed(_T_19) + $signed(_T_20); // @[ChiselImProc.scala 50:13]
  wire [31:0] _T_24 = $signed(io_a_6) * $signed(io_b_6); // @[ChiselImProc.scala 50:24]
  wire [31:0] _T_27 = $signed(_T_23) + $signed(_T_24); // @[ChiselImProc.scala 50:13]
  wire [31:0] _T_28 = $signed(io_a_7) * $signed(io_b_7); // @[ChiselImProc.scala 50:24]
  wire [31:0] _T_31 = $signed(_T_27) + $signed(_T_28); // @[ChiselImProc.scala 50:13]
  wire [31:0] _T_32 = -16'sh1 * $signed(io_b_8); // @[ChiselImProc.scala 50:24]
  assign io_output = $signed(_T_31) + $signed(_T_32); // @[ChiselImProc.scala 53:15]
endmodule
module SqrtExtractionUInt(
  input  [31:0] io_z,
  output [15:0] io_q
);
  wire [32:0] zj_15 = {1'h0,io_z[31:30],30'h0}; // @[Cat.scala 29:58]
  wire [2:0] _T_5 = zj_15[32:30] - 3'h1; // @[Sqrt.scala 54:77]
  wire [32:0] rj_15 = {_T_5,30'h0}; // @[Cat.scala 29:58]
  wire  qSub_15 = ~rj_15[32]; // @[Sqrt.scala 55:27]
  wire [4:0] _T_11 = {rj_15[32:30],io_z[29:28]}; // @[Cat.scala 29:58]
  wire [32:0] _GEN_15 = {_T_11, 28'h0}; // @[Sqrt.scala 59:77]
  wire [35:0] _T_12 = {{3'd0}, _GEN_15}; // @[Sqrt.scala 59:77]
  wire [4:0] _T_15 = {zj_15[32:30],io_z[29:28]}; // @[Cat.scala 29:58]
  wire [32:0] _GEN_16 = {_T_15, 28'h0}; // @[Sqrt.scala 61:77]
  wire [35:0] _T_16 = {{3'd0}, _GEN_16}; // @[Sqrt.scala 61:77]
  wire [35:0] _GEN_0 = qSub_15 ? _T_12 : _T_16; // @[Sqrt.scala 58:26]
  wire [32:0] zj_14 = _GEN_0[32:0]; // @[Sqrt.scala 47:19 Sqrt.scala 59:19 Sqrt.scala 61:19]
  wire [2:0] _T_20 = {qSub_15,2'h1}; // @[Cat.scala 29:58]
  wire [4:0] _GEN_17 = {{2'd0}, _T_20}; // @[Sqrt.scala 64:45]
  wire [4:0] _T_22 = zj_14[32:28] - _GEN_17; // @[Sqrt.scala 64:45]
  wire [32:0] _GEN_18 = {_T_22, 28'h0}; // @[Sqrt.scala 64:77]
  wire [35:0] _T_23 = {{3'd0}, _GEN_18}; // @[Sqrt.scala 64:77]
  wire [32:0] rj_14 = _T_23[32:0]; // @[Sqrt.scala 48:19 Sqrt.scala 64:15]
  wire  qSub_14 = ~rj_14[32]; // @[Sqrt.scala 65:20]
  wire [5:0] _T_28 = {rj_14[31:28],io_z[27:26]}; // @[Cat.scala 29:58]
  wire [31:0] _GEN_19 = {_T_28, 26'h0}; // @[Sqrt.scala 59:77]
  wire [36:0] _T_29 = {{5'd0}, _GEN_19}; // @[Sqrt.scala 59:77]
  wire [5:0] _T_32 = {zj_14[31:28],io_z[27:26]}; // @[Cat.scala 29:58]
  wire [31:0] _GEN_20 = {_T_32, 26'h0}; // @[Sqrt.scala 61:77]
  wire [36:0] _T_33 = {{5'd0}, _GEN_20}; // @[Sqrt.scala 61:77]
  wire [36:0] _GEN_1 = qSub_14 ? _T_29 : _T_33; // @[Sqrt.scala 58:26]
  wire [32:0] zj_13 = _GEN_1[32:0]; // @[Sqrt.scala 47:19 Sqrt.scala 59:19 Sqrt.scala 61:19]
  wire [3:0] _T_38 = {qSub_15,qSub_14,2'h1}; // @[Cat.scala 29:58]
  wire [5:0] _GEN_21 = {{2'd0}, _T_38}; // @[Sqrt.scala 64:45]
  wire [5:0] _T_40 = zj_13[31:26] - _GEN_21; // @[Sqrt.scala 64:45]
  wire [31:0] _GEN_22 = {_T_40, 26'h0}; // @[Sqrt.scala 64:77]
  wire [36:0] _T_41 = {{5'd0}, _GEN_22}; // @[Sqrt.scala 64:77]
  wire [32:0] rj_13 = _T_41[32:0]; // @[Sqrt.scala 48:19 Sqrt.scala 64:15]
  wire  qSub_13 = ~rj_13[31]; // @[Sqrt.scala 65:20]
  wire [6:0] _T_46 = {rj_13[30:26],io_z[25:24]}; // @[Cat.scala 29:58]
  wire [30:0] _GEN_23 = {_T_46, 24'h0}; // @[Sqrt.scala 59:77]
  wire [37:0] _T_47 = {{7'd0}, _GEN_23}; // @[Sqrt.scala 59:77]
  wire [6:0] _T_50 = {zj_13[30:26],io_z[25:24]}; // @[Cat.scala 29:58]
  wire [30:0] _GEN_24 = {_T_50, 24'h0}; // @[Sqrt.scala 61:77]
  wire [37:0] _T_51 = {{7'd0}, _GEN_24}; // @[Sqrt.scala 61:77]
  wire [37:0] _GEN_2 = qSub_13 ? _T_47 : _T_51; // @[Sqrt.scala 58:26]
  wire [32:0] zj_12 = _GEN_2[32:0]; // @[Sqrt.scala 47:19 Sqrt.scala 59:19 Sqrt.scala 61:19]
  wire [4:0] _T_57 = {qSub_15,qSub_14,qSub_13,2'h1}; // @[Cat.scala 29:58]
  wire [6:0] _GEN_25 = {{2'd0}, _T_57}; // @[Sqrt.scala 64:45]
  wire [6:0] _T_59 = zj_12[30:24] - _GEN_25; // @[Sqrt.scala 64:45]
  wire [30:0] _GEN_26 = {_T_59, 24'h0}; // @[Sqrt.scala 64:77]
  wire [37:0] _T_60 = {{7'd0}, _GEN_26}; // @[Sqrt.scala 64:77]
  wire [32:0] rj_12 = _T_60[32:0]; // @[Sqrt.scala 48:19 Sqrt.scala 64:15]
  wire  qSub_12 = ~rj_12[30]; // @[Sqrt.scala 65:20]
  wire [7:0] _T_65 = {rj_12[29:24],io_z[23:22]}; // @[Cat.scala 29:58]
  wire [29:0] _GEN_27 = {_T_65, 22'h0}; // @[Sqrt.scala 59:77]
  wire [38:0] _T_66 = {{9'd0}, _GEN_27}; // @[Sqrt.scala 59:77]
  wire [7:0] _T_69 = {zj_12[29:24],io_z[23:22]}; // @[Cat.scala 29:58]
  wire [29:0] _GEN_28 = {_T_69, 22'h0}; // @[Sqrt.scala 61:77]
  wire [38:0] _T_70 = {{9'd0}, _GEN_28}; // @[Sqrt.scala 61:77]
  wire [38:0] _GEN_3 = qSub_12 ? _T_66 : _T_70; // @[Sqrt.scala 58:26]
  wire [32:0] zj_11 = _GEN_3[32:0]; // @[Sqrt.scala 47:19 Sqrt.scala 59:19 Sqrt.scala 61:19]
  wire [5:0] _T_77 = {qSub_15,qSub_14,qSub_13,qSub_12,2'h1}; // @[Cat.scala 29:58]
  wire [7:0] _GEN_29 = {{2'd0}, _T_77}; // @[Sqrt.scala 64:45]
  wire [7:0] _T_79 = zj_11[29:22] - _GEN_29; // @[Sqrt.scala 64:45]
  wire [29:0] _GEN_30 = {_T_79, 22'h0}; // @[Sqrt.scala 64:77]
  wire [38:0] _T_80 = {{9'd0}, _GEN_30}; // @[Sqrt.scala 64:77]
  wire [32:0] rj_11 = _T_80[32:0]; // @[Sqrt.scala 48:19 Sqrt.scala 64:15]
  wire  qSub_11 = ~rj_11[29]; // @[Sqrt.scala 65:20]
  wire [8:0] _T_85 = {rj_11[28:22],io_z[21:20]}; // @[Cat.scala 29:58]
  wire [28:0] _GEN_31 = {_T_85, 20'h0}; // @[Sqrt.scala 59:77]
  wire [39:0] _T_86 = {{11'd0}, _GEN_31}; // @[Sqrt.scala 59:77]
  wire [8:0] _T_89 = {zj_11[28:22],io_z[21:20]}; // @[Cat.scala 29:58]
  wire [28:0] _GEN_32 = {_T_89, 20'h0}; // @[Sqrt.scala 61:77]
  wire [39:0] _T_90 = {{11'd0}, _GEN_32}; // @[Sqrt.scala 61:77]
  wire [39:0] _GEN_4 = qSub_11 ? _T_86 : _T_90; // @[Sqrt.scala 58:26]
  wire [32:0] zj_10 = _GEN_4[32:0]; // @[Sqrt.scala 47:19 Sqrt.scala 59:19 Sqrt.scala 61:19]
  wire [6:0] _T_98 = {qSub_15,qSub_14,qSub_13,qSub_12,qSub_11,2'h1}; // @[Cat.scala 29:58]
  wire [8:0] _GEN_33 = {{2'd0}, _T_98}; // @[Sqrt.scala 64:45]
  wire [8:0] _T_100 = zj_10[28:20] - _GEN_33; // @[Sqrt.scala 64:45]
  wire [28:0] _GEN_34 = {_T_100, 20'h0}; // @[Sqrt.scala 64:77]
  wire [39:0] _T_101 = {{11'd0}, _GEN_34}; // @[Sqrt.scala 64:77]
  wire [32:0] rj_10 = _T_101[32:0]; // @[Sqrt.scala 48:19 Sqrt.scala 64:15]
  wire  qSub_10 = ~rj_10[28]; // @[Sqrt.scala 65:20]
  wire [9:0] _T_106 = {rj_10[27:20],io_z[19:18]}; // @[Cat.scala 29:58]
  wire [27:0] _GEN_35 = {_T_106, 18'h0}; // @[Sqrt.scala 59:77]
  wire [40:0] _T_107 = {{13'd0}, _GEN_35}; // @[Sqrt.scala 59:77]
  wire [9:0] _T_110 = {zj_10[27:20],io_z[19:18]}; // @[Cat.scala 29:58]
  wire [27:0] _GEN_36 = {_T_110, 18'h0}; // @[Sqrt.scala 61:77]
  wire [40:0] _T_111 = {{13'd0}, _GEN_36}; // @[Sqrt.scala 61:77]
  wire [40:0] _GEN_5 = qSub_10 ? _T_107 : _T_111; // @[Sqrt.scala 58:26]
  wire [32:0] zj_9 = _GEN_5[32:0]; // @[Sqrt.scala 47:19 Sqrt.scala 59:19 Sqrt.scala 61:19]
  wire [7:0] _T_120 = {qSub_15,qSub_14,qSub_13,qSub_12,qSub_11,qSub_10,2'h1}; // @[Cat.scala 29:58]
  wire [9:0] _GEN_37 = {{2'd0}, _T_120}; // @[Sqrt.scala 64:45]
  wire [9:0] _T_122 = zj_9[27:18] - _GEN_37; // @[Sqrt.scala 64:45]
  wire [27:0] _GEN_38 = {_T_122, 18'h0}; // @[Sqrt.scala 64:77]
  wire [40:0] _T_123 = {{13'd0}, _GEN_38}; // @[Sqrt.scala 64:77]
  wire [32:0] rj_9 = _T_123[32:0]; // @[Sqrt.scala 48:19 Sqrt.scala 64:15]
  wire  qSub_9 = ~rj_9[27]; // @[Sqrt.scala 65:20]
  wire [10:0] _T_128 = {rj_9[26:18],io_z[17:16]}; // @[Cat.scala 29:58]
  wire [26:0] _GEN_39 = {_T_128, 16'h0}; // @[Sqrt.scala 59:77]
  wire [41:0] _T_129 = {{15'd0}, _GEN_39}; // @[Sqrt.scala 59:77]
  wire [10:0] _T_132 = {zj_9[26:18],io_z[17:16]}; // @[Cat.scala 29:58]
  wire [26:0] _GEN_40 = {_T_132, 16'h0}; // @[Sqrt.scala 61:77]
  wire [41:0] _T_133 = {{15'd0}, _GEN_40}; // @[Sqrt.scala 61:77]
  wire [41:0] _GEN_6 = qSub_9 ? _T_129 : _T_133; // @[Sqrt.scala 58:26]
  wire [32:0] zj_8 = _GEN_6[32:0]; // @[Sqrt.scala 47:19 Sqrt.scala 59:19 Sqrt.scala 61:19]
  wire [8:0] _T_143 = {qSub_15,qSub_14,qSub_13,qSub_12,qSub_11,qSub_10,qSub_9,2'h1}; // @[Cat.scala 29:58]
  wire [10:0] _GEN_41 = {{2'd0}, _T_143}; // @[Sqrt.scala 64:45]
  wire [10:0] _T_145 = zj_8[26:16] - _GEN_41; // @[Sqrt.scala 64:45]
  wire [26:0] _GEN_42 = {_T_145, 16'h0}; // @[Sqrt.scala 64:77]
  wire [41:0] _T_146 = {{15'd0}, _GEN_42}; // @[Sqrt.scala 64:77]
  wire [32:0] rj_8 = _T_146[32:0]; // @[Sqrt.scala 48:19 Sqrt.scala 64:15]
  wire  qSub_8 = ~rj_8[26]; // @[Sqrt.scala 65:20]
  wire [11:0] _T_151 = {rj_8[25:16],io_z[15:14]}; // @[Cat.scala 29:58]
  wire [25:0] _GEN_43 = {_T_151, 14'h0}; // @[Sqrt.scala 59:77]
  wire [26:0] _T_152 = {{1'd0}, _GEN_43}; // @[Sqrt.scala 59:77]
  wire [11:0] _T_155 = {zj_8[25:16],io_z[15:14]}; // @[Cat.scala 29:58]
  wire [25:0] _GEN_44 = {_T_155, 14'h0}; // @[Sqrt.scala 61:77]
  wire [26:0] _T_156 = {{1'd0}, _GEN_44}; // @[Sqrt.scala 61:77]
  wire [26:0] _GEN_7 = qSub_8 ? _T_152 : _T_156; // @[Sqrt.scala 58:26]
  wire [32:0] zj_7 = {{6'd0}, _GEN_7}; // @[Sqrt.scala 47:19 Sqrt.scala 59:19 Sqrt.scala 61:19]
  wire [7:0] _T_166 = {qSub_15,qSub_14,qSub_13,qSub_12,qSub_11,qSub_10,qSub_9,qSub_8}; // @[Sqrt.scala 64:58]
  wire [9:0] _T_167 = {qSub_15,qSub_14,qSub_13,qSub_12,qSub_11,qSub_10,qSub_9,qSub_8,2'h1}; // @[Cat.scala 29:58]
  wire [11:0] _GEN_45 = {{2'd0}, _T_167}; // @[Sqrt.scala 64:45]
  wire [11:0] _T_169 = zj_7[25:14] - _GEN_45; // @[Sqrt.scala 64:45]
  wire [25:0] _GEN_46 = {_T_169, 14'h0}; // @[Sqrt.scala 64:77]
  wire [26:0] _T_170 = {{1'd0}, _GEN_46}; // @[Sqrt.scala 64:77]
  wire [32:0] rj_7 = {{6'd0}, _T_170}; // @[Sqrt.scala 48:19 Sqrt.scala 64:15]
  wire  qSub_7 = ~rj_7[25]; // @[Sqrt.scala 65:20]
  wire [12:0] _T_175 = {rj_7[24:14],io_z[13:12]}; // @[Cat.scala 29:58]
  wire [24:0] _GEN_47 = {_T_175, 12'h0}; // @[Sqrt.scala 59:77]
  wire [27:0] _T_176 = {{3'd0}, _GEN_47}; // @[Sqrt.scala 59:77]
  wire [12:0] _T_179 = {zj_7[24:14],io_z[13:12]}; // @[Cat.scala 29:58]
  wire [24:0] _GEN_48 = {_T_179, 12'h0}; // @[Sqrt.scala 61:77]
  wire [27:0] _T_180 = {{3'd0}, _GEN_48}; // @[Sqrt.scala 61:77]
  wire [27:0] _GEN_8 = qSub_7 ? _T_176 : _T_180; // @[Sqrt.scala 58:26]
  wire [32:0] zj_6 = {{5'd0}, _GEN_8}; // @[Sqrt.scala 47:19 Sqrt.scala 59:19 Sqrt.scala 61:19]
  wire [10:0] _T_192 = {qSub_15,qSub_14,qSub_13,qSub_12,qSub_11,qSub_10,qSub_9,qSub_8,qSub_7,2'h1}; // @[Cat.scala 29:58]
  wire [12:0] _GEN_49 = {{2'd0}, _T_192}; // @[Sqrt.scala 64:45]
  wire [12:0] _T_194 = zj_6[24:12] - _GEN_49; // @[Sqrt.scala 64:45]
  wire [24:0] _GEN_50 = {_T_194, 12'h0}; // @[Sqrt.scala 64:77]
  wire [27:0] _T_195 = {{3'd0}, _GEN_50}; // @[Sqrt.scala 64:77]
  wire [32:0] rj_6 = {{5'd0}, _T_195}; // @[Sqrt.scala 48:19 Sqrt.scala 64:15]
  wire  qSub_6 = ~rj_6[24]; // @[Sqrt.scala 65:20]
  wire [13:0] _T_200 = {rj_6[23:12],io_z[11:10]}; // @[Cat.scala 29:58]
  wire [23:0] _GEN_51 = {_T_200, 10'h0}; // @[Sqrt.scala 59:77]
  wire [28:0] _T_201 = {{5'd0}, _GEN_51}; // @[Sqrt.scala 59:77]
  wire [13:0] _T_204 = {zj_6[23:12],io_z[11:10]}; // @[Cat.scala 29:58]
  wire [23:0] _GEN_52 = {_T_204, 10'h0}; // @[Sqrt.scala 61:77]
  wire [28:0] _T_205 = {{5'd0}, _GEN_52}; // @[Sqrt.scala 61:77]
  wire [28:0] _GEN_9 = qSub_6 ? _T_201 : _T_205; // @[Sqrt.scala 58:26]
  wire [32:0] zj_5 = {{4'd0}, _GEN_9}; // @[Sqrt.scala 47:19 Sqrt.scala 59:19 Sqrt.scala 61:19]
  wire [9:0] _T_217 = {qSub_15,qSub_14,qSub_13,qSub_12,qSub_11,qSub_10,qSub_9,qSub_8,qSub_7,qSub_6}; // @[Sqrt.scala 64:58]
  wire [11:0] _T_218 = {_T_217,2'h1}; // @[Cat.scala 29:58]
  wire [13:0] _GEN_53 = {{2'd0}, _T_218}; // @[Sqrt.scala 64:45]
  wire [13:0] _T_220 = zj_5[23:10] - _GEN_53; // @[Sqrt.scala 64:45]
  wire [23:0] _GEN_54 = {_T_220, 10'h0}; // @[Sqrt.scala 64:77]
  wire [28:0] _T_221 = {{5'd0}, _GEN_54}; // @[Sqrt.scala 64:77]
  wire [32:0] rj_5 = {{4'd0}, _T_221}; // @[Sqrt.scala 48:19 Sqrt.scala 64:15]
  wire  qSub_5 = ~rj_5[23]; // @[Sqrt.scala 65:20]
  wire [14:0] _T_226 = {rj_5[22:10],io_z[9:8]}; // @[Cat.scala 29:58]
  wire [22:0] _GEN_55 = {_T_226, 8'h0}; // @[Sqrt.scala 59:77]
  wire [29:0] _T_227 = {{7'd0}, _GEN_55}; // @[Sqrt.scala 59:77]
  wire [14:0] _T_230 = {zj_5[22:10],io_z[9:8]}; // @[Cat.scala 29:58]
  wire [22:0] _GEN_56 = {_T_230, 8'h0}; // @[Sqrt.scala 61:77]
  wire [29:0] _T_231 = {{7'd0}, _GEN_56}; // @[Sqrt.scala 61:77]
  wire [29:0] _GEN_10 = qSub_5 ? _T_227 : _T_231; // @[Sqrt.scala 58:26]
  wire [32:0] zj_4 = {{3'd0}, _GEN_10}; // @[Sqrt.scala 47:19 Sqrt.scala 59:19 Sqrt.scala 61:19]
  wire [4:0] _T_238 = {qSub_9,qSub_8,qSub_7,qSub_6,qSub_5}; // @[Sqrt.scala 64:58]
  wire [12:0] _T_245 = {qSub_15,qSub_14,qSub_13,qSub_12,qSub_11,qSub_10,_T_238,2'h1}; // @[Cat.scala 29:58]
  wire [14:0] _GEN_57 = {{2'd0}, _T_245}; // @[Sqrt.scala 64:45]
  wire [14:0] _T_247 = zj_4[22:8] - _GEN_57; // @[Sqrt.scala 64:45]
  wire [22:0] _GEN_58 = {_T_247, 8'h0}; // @[Sqrt.scala 64:77]
  wire [29:0] _T_248 = {{7'd0}, _GEN_58}; // @[Sqrt.scala 64:77]
  wire [32:0] rj_4 = {{3'd0}, _T_248}; // @[Sqrt.scala 48:19 Sqrt.scala 64:15]
  wire  qSub_4 = ~rj_4[22]; // @[Sqrt.scala 65:20]
  wire [15:0] _T_253 = {rj_4[21:8],io_z[7:6]}; // @[Cat.scala 29:58]
  wire [21:0] _GEN_59 = {_T_253, 6'h0}; // @[Sqrt.scala 59:77]
  wire [22:0] _T_254 = {{1'd0}, _GEN_59}; // @[Sqrt.scala 59:77]
  wire [15:0] _T_257 = {zj_4[21:8],io_z[7:6]}; // @[Cat.scala 29:58]
  wire [21:0] _GEN_60 = {_T_257, 6'h0}; // @[Sqrt.scala 61:77]
  wire [22:0] _T_258 = {{1'd0}, _GEN_60}; // @[Sqrt.scala 61:77]
  wire [22:0] _GEN_11 = qSub_4 ? _T_254 : _T_258; // @[Sqrt.scala 58:26]
  wire [32:0] zj_3 = {{10'd0}, _GEN_11}; // @[Sqrt.scala 47:19 Sqrt.scala 59:19 Sqrt.scala 61:19]
  wire [5:0] _T_266 = {qSub_9,qSub_8,qSub_7,qSub_6,qSub_5,qSub_4}; // @[Sqrt.scala 64:58]
  wire [13:0] _T_273 = {qSub_15,qSub_14,qSub_13,qSub_12,qSub_11,qSub_10,_T_266,2'h1}; // @[Cat.scala 29:58]
  wire [15:0] _GEN_61 = {{2'd0}, _T_273}; // @[Sqrt.scala 64:45]
  wire [15:0] _T_275 = zj_3[21:6] - _GEN_61; // @[Sqrt.scala 64:45]
  wire [21:0] _GEN_62 = {_T_275, 6'h0}; // @[Sqrt.scala 64:77]
  wire [22:0] _T_276 = {{1'd0}, _GEN_62}; // @[Sqrt.scala 64:77]
  wire [32:0] rj_3 = {{10'd0}, _T_276}; // @[Sqrt.scala 48:19 Sqrt.scala 64:15]
  wire  qSub_3 = ~rj_3[21]; // @[Sqrt.scala 65:20]
  wire [16:0] _T_281 = {rj_3[20:6],io_z[5:4]}; // @[Cat.scala 29:58]
  wire [20:0] _GEN_63 = {_T_281, 4'h0}; // @[Sqrt.scala 59:77]
  wire [23:0] _T_282 = {{3'd0}, _GEN_63}; // @[Sqrt.scala 59:77]
  wire [16:0] _T_285 = {zj_3[20:6],io_z[5:4]}; // @[Cat.scala 29:58]
  wire [20:0] _GEN_64 = {_T_285, 4'h0}; // @[Sqrt.scala 61:77]
  wire [23:0] _T_286 = {{3'd0}, _GEN_64}; // @[Sqrt.scala 61:77]
  wire [23:0] _GEN_12 = qSub_3 ? _T_282 : _T_286; // @[Sqrt.scala 58:26]
  wire [32:0] zj_2 = {{9'd0}, _GEN_12}; // @[Sqrt.scala 47:19 Sqrt.scala 59:19 Sqrt.scala 61:19]
  wire [5:0] _T_294 = {qSub_8,qSub_7,qSub_6,qSub_5,qSub_4,qSub_3}; // @[Sqrt.scala 64:58]
  wire [14:0] _T_302 = {qSub_15,qSub_14,qSub_13,qSub_12,qSub_11,qSub_10,qSub_9,_T_294,2'h1}; // @[Cat.scala 29:58]
  wire [16:0] _GEN_65 = {{2'd0}, _T_302}; // @[Sqrt.scala 64:45]
  wire [16:0] _T_304 = zj_2[20:4] - _GEN_65; // @[Sqrt.scala 64:45]
  wire [20:0] _GEN_66 = {_T_304, 4'h0}; // @[Sqrt.scala 64:77]
  wire [23:0] _T_305 = {{3'd0}, _GEN_66}; // @[Sqrt.scala 64:77]
  wire [32:0] rj_2 = {{9'd0}, _T_305}; // @[Sqrt.scala 48:19 Sqrt.scala 64:15]
  wire  qSub_2 = ~rj_2[20]; // @[Sqrt.scala 65:20]
  wire [17:0] _T_310 = {rj_2[19:4],io_z[3:2]}; // @[Cat.scala 29:58]
  wire [19:0] _GEN_67 = {_T_310, 2'h0}; // @[Sqrt.scala 59:77]
  wire [20:0] _T_311 = {{1'd0}, _GEN_67}; // @[Sqrt.scala 59:77]
  wire [17:0] _T_314 = {zj_2[19:4],io_z[3:2]}; // @[Cat.scala 29:58]
  wire [19:0] _GEN_68 = {_T_314, 2'h0}; // @[Sqrt.scala 61:77]
  wire [20:0] _T_315 = {{1'd0}, _GEN_68}; // @[Sqrt.scala 61:77]
  wire [20:0] _GEN_13 = qSub_2 ? _T_311 : _T_315; // @[Sqrt.scala 58:26]
  wire [32:0] zj_1 = {{12'd0}, _GEN_13}; // @[Sqrt.scala 47:19 Sqrt.scala 59:19 Sqrt.scala 61:19]
  wire [6:0] _T_324 = {qSub_8,qSub_7,qSub_6,qSub_5,qSub_4,qSub_3,qSub_2}; // @[Sqrt.scala 64:58]
  wire [15:0] _T_332 = {qSub_15,qSub_14,qSub_13,qSub_12,qSub_11,qSub_10,qSub_9,_T_324,2'h1}; // @[Cat.scala 29:58]
  wire [17:0] _GEN_69 = {{2'd0}, _T_332}; // @[Sqrt.scala 64:45]
  wire [17:0] _T_334 = zj_1[19:2] - _GEN_69; // @[Sqrt.scala 64:45]
  wire [19:0] _GEN_70 = {_T_334, 2'h0}; // @[Sqrt.scala 64:77]
  wire [20:0] _T_335 = {{1'd0}, _GEN_70}; // @[Sqrt.scala 64:77]
  wire [32:0] rj_1 = {{12'd0}, _T_335}; // @[Sqrt.scala 48:19 Sqrt.scala 64:15]
  wire  qSub_1 = ~rj_1[19]; // @[Sqrt.scala 65:20]
  wire [18:0] _T_340 = {rj_1[18:2],io_z[1:0]}; // @[Cat.scala 29:58]
  wire [19:0] _T_341 = {{1'd0}, _T_340}; // @[Sqrt.scala 59:77]
  wire [18:0] _T_344 = {zj_1[18:2],io_z[1:0]}; // @[Cat.scala 29:58]
  wire [19:0] _T_345 = {{1'd0}, _T_344}; // @[Sqrt.scala 61:77]
  wire [19:0] _GEN_14 = qSub_1 ? _T_341 : _T_345; // @[Sqrt.scala 58:26]
  wire [32:0] zj_0 = {{13'd0}, _GEN_14}; // @[Sqrt.scala 47:19 Sqrt.scala 59:19 Sqrt.scala 61:19]
  wire [6:0] _T_354 = {qSub_7,qSub_6,qSub_5,qSub_4,qSub_3,qSub_2,qSub_1}; // @[Sqrt.scala 64:58]
  wire [16:0] _T_363 = {qSub_15,qSub_14,qSub_13,qSub_12,qSub_11,qSub_10,qSub_9,qSub_8,_T_354,2'h1}; // @[Cat.scala 29:58]
  wire [18:0] _GEN_71 = {{2'd0}, _T_363}; // @[Sqrt.scala 64:45]
  wire [18:0] _T_365 = zj_0[18:0] - _GEN_71; // @[Sqrt.scala 64:45]
  wire [19:0] _T_366 = {{1'd0}, _T_365}; // @[Sqrt.scala 64:77]
  wire [32:0] rj_0 = {{13'd0}, _T_366}; // @[Sqrt.scala 48:19 Sqrt.scala 64:15]
  wire  qSub_0 = ~rj_0[18]; // @[Sqrt.scala 65:20]
  wire [7:0] _T_375 = {qSub_7,qSub_6,qSub_5,qSub_4,qSub_3,qSub_2,qSub_1,qSub_0}; // @[Sqrt.scala 68:18]
  assign io_q = {_T_166,_T_375}; // @[Sqrt.scala 68:10]
endmodule
module SobelFilter(
  input        clock,
  input        reset,
  output       io_enq_ready,
  input        io_enq_valid,
  input  [7:0] io_enq_bits,
  input        io_enq_user,
  input        io_enq_last,
  input        io_deq_ready,
  output       io_deq_valid,
  output [1:0] io_deq_bits_grad_dir,
  output [7:0] io_deq_bits_value,
  output       io_deq_user,
  output       io_deq_last
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
  reg [31:0] _RAND_64;
  reg [31:0] _RAND_65;
  reg [31:0] _RAND_66;
  reg [31:0] _RAND_67;
  reg [31:0] _RAND_68;
  reg [31:0] _RAND_69;
  reg [31:0] _RAND_70;
  reg [31:0] _RAND_71;
  reg [31:0] _RAND_72;
  reg [31:0] _RAND_73;
  reg [31:0] _RAND_74;
  reg [31:0] _RAND_75;
  reg [31:0] _RAND_76;
  reg [31:0] _RAND_77;
  reg [31:0] _RAND_78;
  reg [31:0] _RAND_79;
  reg [31:0] _RAND_80;
  reg [31:0] _RAND_81;
  reg [31:0] _RAND_82;
  reg [31:0] _RAND_83;
  reg [31:0] _RAND_84;
  reg [31:0] _RAND_85;
  reg [31:0] _RAND_86;
  reg [31:0] _RAND_87;
  reg [31:0] _RAND_88;
  reg [31:0] _RAND_89;
  reg [31:0] _RAND_90;
  reg [31:0] _RAND_91;
  reg [31:0] _RAND_92;
  reg [31:0] _RAND_93;
  reg [31:0] _RAND_94;
  reg [31:0] _RAND_95;
  reg [31:0] _RAND_96;
  reg [31:0] _RAND_97;
  reg [31:0] _RAND_98;
  reg [31:0] _RAND_99;
  reg [31:0] _RAND_100;
  reg [31:0] _RAND_101;
  reg [31:0] _RAND_102;
  reg [31:0] _RAND_103;
  reg [31:0] _RAND_104;
  reg [31:0] _RAND_105;
  reg [31:0] _RAND_106;
  reg [31:0] _RAND_107;
  reg [31:0] _RAND_108;
  reg [31:0] _RAND_109;
  reg [31:0] _RAND_110;
  reg [31:0] _RAND_111;
  reg [31:0] _RAND_112;
  reg [31:0] _RAND_113;
  reg [31:0] _RAND_114;
  reg [31:0] _RAND_115;
  reg [31:0] _RAND_116;
  reg [31:0] _RAND_117;
  reg [31:0] _RAND_118;
  reg [31:0] _RAND_119;
  reg [31:0] _RAND_120;
  reg [31:0] _RAND_121;
  reg [31:0] _RAND_122;
  reg [31:0] _RAND_123;
  reg [31:0] _RAND_124;
  reg [31:0] _RAND_125;
  reg [31:0] _RAND_126;
  reg [31:0] _RAND_127;
  reg [31:0] _RAND_128;
  reg [31:0] _RAND_129;
  reg [31:0] _RAND_130;
  reg [31:0] _RAND_131;
  reg [31:0] _RAND_132;
  reg [31:0] _RAND_133;
  reg [31:0] _RAND_134;
  reg [31:0] _RAND_135;
  reg [31:0] _RAND_136;
  reg [31:0] _RAND_137;
  reg [31:0] _RAND_138;
  reg [31:0] _RAND_139;
  reg [31:0] _RAND_140;
  reg [31:0] _RAND_141;
  reg [31:0] _RAND_142;
  reg [31:0] _RAND_143;
  reg [31:0] _RAND_144;
  reg [31:0] _RAND_145;
  reg [31:0] _RAND_146;
  reg [31:0] _RAND_147;
  reg [31:0] _RAND_148;
  reg [31:0] _RAND_149;
  reg [31:0] _RAND_150;
  reg [31:0] _RAND_151;
  reg [31:0] _RAND_152;
  reg [31:0] _RAND_153;
  reg [31:0] _RAND_154;
  reg [31:0] _RAND_155;
  reg [31:0] _RAND_156;
  reg [31:0] _RAND_157;
  reg [31:0] _RAND_158;
  reg [31:0] _RAND_159;
  reg [31:0] _RAND_160;
  reg [31:0] _RAND_161;
  reg [31:0] _RAND_162;
  reg [31:0] _RAND_163;
  reg [31:0] _RAND_164;
  reg [31:0] _RAND_165;
  reg [31:0] _RAND_166;
  reg [31:0] _RAND_167;
  reg [31:0] _RAND_168;
  reg [31:0] _RAND_169;
  reg [31:0] _RAND_170;
  reg [31:0] _RAND_171;
  reg [31:0] _RAND_172;
  reg [31:0] _RAND_173;
  reg [31:0] _RAND_174;
  reg [31:0] _RAND_175;
  reg [31:0] _RAND_176;
  reg [31:0] _RAND_177;
  reg [31:0] _RAND_178;
  reg [31:0] _RAND_179;
  reg [31:0] _RAND_180;
  reg [31:0] _RAND_181;
  reg [31:0] _RAND_182;
  reg [31:0] _RAND_183;
  reg [31:0] _RAND_184;
  reg [31:0] _RAND_185;
  reg [31:0] _RAND_186;
  reg [31:0] _RAND_187;
  reg [31:0] _RAND_188;
  reg [31:0] _RAND_189;
  reg [31:0] _RAND_190;
  reg [31:0] _RAND_191;
  reg [31:0] _RAND_192;
  reg [31:0] _RAND_193;
  reg [31:0] _RAND_194;
  reg [31:0] _RAND_195;
  reg [31:0] _RAND_196;
  reg [31:0] _RAND_197;
  reg [31:0] _RAND_198;
  reg [31:0] _RAND_199;
  reg [31:0] _RAND_200;
  reg [31:0] _RAND_201;
  reg [31:0] _RAND_202;
  reg [31:0] _RAND_203;
  reg [31:0] _RAND_204;
  reg [31:0] _RAND_205;
  reg [31:0] _RAND_206;
  reg [31:0] _RAND_207;
  reg [31:0] _RAND_208;
  reg [31:0] _RAND_209;
  reg [31:0] _RAND_210;
  reg [31:0] _RAND_211;
  reg [31:0] _RAND_212;
  reg [31:0] _RAND_213;
  reg [31:0] _RAND_214;
  reg [31:0] _RAND_215;
  reg [31:0] _RAND_216;
  reg [31:0] _RAND_217;
  reg [31:0] _RAND_218;
  reg [31:0] _RAND_219;
  reg [31:0] _RAND_220;
  reg [31:0] _RAND_221;
  reg [31:0] _RAND_222;
  reg [31:0] _RAND_223;
  reg [31:0] _RAND_224;
  reg [31:0] _RAND_225;
  reg [31:0] _RAND_226;
  reg [31:0] _RAND_227;
  reg [31:0] _RAND_228;
  reg [31:0] _RAND_229;
  reg [31:0] _RAND_230;
  reg [31:0] _RAND_231;
  reg [31:0] _RAND_232;
  reg [31:0] _RAND_233;
  reg [31:0] _RAND_234;
  reg [31:0] _RAND_235;
  reg [31:0] _RAND_236;
  reg [31:0] _RAND_237;
  reg [31:0] _RAND_238;
  reg [31:0] _RAND_239;
  reg [31:0] _RAND_240;
  reg [31:0] _RAND_241;
  reg [31:0] _RAND_242;
  reg [31:0] _RAND_243;
  reg [31:0] _RAND_244;
  reg [31:0] _RAND_245;
  reg [31:0] _RAND_246;
  reg [31:0] _RAND_247;
  reg [31:0] _RAND_248;
  reg [31:0] _RAND_249;
  reg [31:0] _RAND_250;
  reg [31:0] _RAND_251;
  reg [31:0] _RAND_252;
  reg [31:0] _RAND_253;
  reg [31:0] _RAND_254;
  reg [31:0] _RAND_255;
  reg [31:0] _RAND_256;
  reg [31:0] _RAND_257;
  reg [31:0] _RAND_258;
  reg [31:0] _RAND_259;
  reg [31:0] _RAND_260;
  reg [31:0] _RAND_261;
  reg [31:0] _RAND_262;
  reg [31:0] _RAND_263;
  reg [31:0] _RAND_264;
  reg [31:0] _RAND_265;
  reg [31:0] _RAND_266;
  reg [31:0] _RAND_267;
  reg [31:0] _RAND_268;
  reg [31:0] _RAND_269;
  reg [31:0] _RAND_270;
  reg [31:0] _RAND_271;
  reg [31:0] _RAND_272;
  reg [31:0] _RAND_273;
  reg [31:0] _RAND_274;
  reg [31:0] _RAND_275;
  reg [31:0] _RAND_276;
  reg [31:0] _RAND_277;
  reg [31:0] _RAND_278;
  reg [31:0] _RAND_279;
  reg [31:0] _RAND_280;
  reg [31:0] _RAND_281;
  reg [31:0] _RAND_282;
  reg [31:0] _RAND_283;
  reg [31:0] _RAND_284;
  reg [31:0] _RAND_285;
  reg [31:0] _RAND_286;
  reg [31:0] _RAND_287;
  reg [31:0] _RAND_288;
  reg [31:0] _RAND_289;
  reg [31:0] _RAND_290;
  reg [31:0] _RAND_291;
  reg [31:0] _RAND_292;
  reg [31:0] _RAND_293;
  reg [31:0] _RAND_294;
  reg [31:0] _RAND_295;
  reg [31:0] _RAND_296;
  reg [31:0] _RAND_297;
  reg [31:0] _RAND_298;
  reg [31:0] _RAND_299;
  reg [31:0] _RAND_300;
  reg [31:0] _RAND_301;
  reg [31:0] _RAND_302;
  reg [31:0] _RAND_303;
  reg [31:0] _RAND_304;
  reg [31:0] _RAND_305;
  reg [31:0] _RAND_306;
  reg [31:0] _RAND_307;
  reg [31:0] _RAND_308;
  reg [31:0] _RAND_309;
  reg [31:0] _RAND_310;
  reg [31:0] _RAND_311;
  reg [31:0] _RAND_312;
  reg [31:0] _RAND_313;
  reg [31:0] _RAND_314;
  reg [31:0] _RAND_315;
  reg [31:0] _RAND_316;
  reg [31:0] _RAND_317;
  reg [31:0] _RAND_318;
  reg [31:0] _RAND_319;
  reg [31:0] _RAND_320;
  reg [31:0] _RAND_321;
  reg [31:0] _RAND_322;
  reg [31:0] _RAND_323;
  reg [31:0] _RAND_324;
  reg [31:0] _RAND_325;
  reg [31:0] _RAND_326;
  reg [31:0] _RAND_327;
  reg [31:0] _RAND_328;
  reg [31:0] _RAND_329;
  reg [31:0] _RAND_330;
  reg [31:0] _RAND_331;
  reg [31:0] _RAND_332;
  reg [31:0] _RAND_333;
  reg [31:0] _RAND_334;
  reg [31:0] _RAND_335;
  reg [31:0] _RAND_336;
  reg [31:0] _RAND_337;
  reg [31:0] _RAND_338;
  reg [31:0] _RAND_339;
  reg [31:0] _RAND_340;
  reg [31:0] _RAND_341;
  reg [31:0] _RAND_342;
  reg [31:0] _RAND_343;
  reg [31:0] _RAND_344;
  reg [31:0] _RAND_345;
  reg [31:0] _RAND_346;
  reg [31:0] _RAND_347;
  reg [31:0] _RAND_348;
  reg [31:0] _RAND_349;
  reg [31:0] _RAND_350;
  reg [31:0] _RAND_351;
  reg [31:0] _RAND_352;
  reg [31:0] _RAND_353;
  reg [31:0] _RAND_354;
  reg [31:0] _RAND_355;
  reg [31:0] _RAND_356;
  reg [31:0] _RAND_357;
  reg [31:0] _RAND_358;
  reg [31:0] _RAND_359;
  reg [31:0] _RAND_360;
  reg [31:0] _RAND_361;
  reg [31:0] _RAND_362;
  reg [31:0] _RAND_363;
  reg [31:0] _RAND_364;
  reg [31:0] _RAND_365;
  reg [31:0] _RAND_366;
  reg [31:0] _RAND_367;
  reg [31:0] _RAND_368;
  reg [31:0] _RAND_369;
  reg [31:0] _RAND_370;
  reg [31:0] _RAND_371;
  reg [31:0] _RAND_372;
  reg [31:0] _RAND_373;
  reg [31:0] _RAND_374;
  reg [31:0] _RAND_375;
  reg [31:0] _RAND_376;
  reg [31:0] _RAND_377;
  reg [31:0] _RAND_378;
  reg [31:0] _RAND_379;
  reg [31:0] _RAND_380;
  reg [31:0] _RAND_381;
  reg [31:0] _RAND_382;
  reg [31:0] _RAND_383;
  reg [31:0] _RAND_384;
  reg [31:0] _RAND_385;
  reg [31:0] _RAND_386;
  reg [31:0] _RAND_387;
  reg [31:0] _RAND_388;
  reg [31:0] _RAND_389;
  reg [31:0] _RAND_390;
  reg [31:0] _RAND_391;
  reg [31:0] _RAND_392;
  reg [31:0] _RAND_393;
  reg [31:0] _RAND_394;
  reg [31:0] _RAND_395;
  reg [31:0] _RAND_396;
  reg [31:0] _RAND_397;
  reg [31:0] _RAND_398;
  reg [31:0] _RAND_399;
  reg [31:0] _RAND_400;
  reg [31:0] _RAND_401;
  reg [31:0] _RAND_402;
  reg [31:0] _RAND_403;
  reg [31:0] _RAND_404;
  reg [31:0] _RAND_405;
  reg [31:0] _RAND_406;
  reg [31:0] _RAND_407;
  reg [31:0] _RAND_408;
  reg [31:0] _RAND_409;
  reg [31:0] _RAND_410;
  reg [31:0] _RAND_411;
  reg [31:0] _RAND_412;
  reg [31:0] _RAND_413;
  reg [31:0] _RAND_414;
  reg [31:0] _RAND_415;
  reg [31:0] _RAND_416;
  reg [31:0] _RAND_417;
  reg [31:0] _RAND_418;
  reg [31:0] _RAND_419;
  reg [31:0] _RAND_420;
  reg [31:0] _RAND_421;
  reg [31:0] _RAND_422;
  reg [31:0] _RAND_423;
  reg [31:0] _RAND_424;
  reg [31:0] _RAND_425;
  reg [31:0] _RAND_426;
  reg [31:0] _RAND_427;
  reg [31:0] _RAND_428;
  reg [31:0] _RAND_429;
  reg [31:0] _RAND_430;
  reg [31:0] _RAND_431;
  reg [31:0] _RAND_432;
  reg [31:0] _RAND_433;
  reg [31:0] _RAND_434;
  reg [31:0] _RAND_435;
  reg [31:0] _RAND_436;
  reg [31:0] _RAND_437;
  reg [31:0] _RAND_438;
  reg [31:0] _RAND_439;
  reg [31:0] _RAND_440;
  reg [31:0] _RAND_441;
  reg [31:0] _RAND_442;
  reg [31:0] _RAND_443;
  reg [31:0] _RAND_444;
  reg [31:0] _RAND_445;
  reg [31:0] _RAND_446;
  reg [31:0] _RAND_447;
  reg [31:0] _RAND_448;
  reg [31:0] _RAND_449;
  reg [31:0] _RAND_450;
  reg [31:0] _RAND_451;
  reg [31:0] _RAND_452;
  reg [31:0] _RAND_453;
  reg [31:0] _RAND_454;
  reg [31:0] _RAND_455;
  reg [31:0] _RAND_456;
  reg [31:0] _RAND_457;
  reg [31:0] _RAND_458;
  reg [31:0] _RAND_459;
  reg [31:0] _RAND_460;
  reg [31:0] _RAND_461;
  reg [31:0] _RAND_462;
  reg [31:0] _RAND_463;
  reg [31:0] _RAND_464;
  reg [31:0] _RAND_465;
  reg [31:0] _RAND_466;
  reg [31:0] _RAND_467;
  reg [31:0] _RAND_468;
  reg [31:0] _RAND_469;
  reg [31:0] _RAND_470;
  reg [31:0] _RAND_471;
  reg [31:0] _RAND_472;
  reg [31:0] _RAND_473;
  reg [31:0] _RAND_474;
  reg [31:0] _RAND_475;
  reg [31:0] _RAND_476;
  reg [31:0] _RAND_477;
  reg [31:0] _RAND_478;
  reg [31:0] _RAND_479;
  reg [31:0] _RAND_480;
  reg [31:0] _RAND_481;
  reg [31:0] _RAND_482;
  reg [31:0] _RAND_483;
  reg [31:0] _RAND_484;
  reg [31:0] _RAND_485;
  reg [31:0] _RAND_486;
  reg [31:0] _RAND_487;
  reg [31:0] _RAND_488;
  reg [31:0] _RAND_489;
  reg [31:0] _RAND_490;
  reg [31:0] _RAND_491;
  reg [31:0] _RAND_492;
  reg [31:0] _RAND_493;
  reg [31:0] _RAND_494;
  reg [31:0] _RAND_495;
  reg [31:0] _RAND_496;
  reg [31:0] _RAND_497;
  reg [31:0] _RAND_498;
  reg [31:0] _RAND_499;
  reg [31:0] _RAND_500;
  reg [31:0] _RAND_501;
  reg [31:0] _RAND_502;
  reg [31:0] _RAND_503;
  reg [31:0] _RAND_504;
  reg [31:0] _RAND_505;
  reg [31:0] _RAND_506;
  reg [31:0] _RAND_507;
  reg [31:0] _RAND_508;
  reg [31:0] _RAND_509;
  reg [31:0] _RAND_510;
  reg [31:0] _RAND_511;
  reg [31:0] _RAND_512;
  reg [31:0] _RAND_513;
  reg [31:0] _RAND_514;
  reg [31:0] _RAND_515;
  reg [31:0] _RAND_516;
  reg [31:0] _RAND_517;
  reg [31:0] _RAND_518;
  reg [31:0] _RAND_519;
  reg [31:0] _RAND_520;
  reg [31:0] _RAND_521;
  reg [31:0] _RAND_522;
  reg [31:0] _RAND_523;
  reg [31:0] _RAND_524;
  reg [31:0] _RAND_525;
  reg [31:0] _RAND_526;
  reg [31:0] _RAND_527;
  reg [31:0] _RAND_528;
  reg [31:0] _RAND_529;
  reg [31:0] _RAND_530;
  reg [31:0] _RAND_531;
  reg [31:0] _RAND_532;
  reg [31:0] _RAND_533;
  reg [31:0] _RAND_534;
  reg [31:0] _RAND_535;
  reg [31:0] _RAND_536;
  reg [31:0] _RAND_537;
  reg [31:0] _RAND_538;
  reg [31:0] _RAND_539;
  reg [31:0] _RAND_540;
  reg [31:0] _RAND_541;
  reg [31:0] _RAND_542;
  reg [31:0] _RAND_543;
  reg [31:0] _RAND_544;
  reg [31:0] _RAND_545;
  reg [31:0] _RAND_546;
  reg [31:0] _RAND_547;
  reg [31:0] _RAND_548;
  reg [31:0] _RAND_549;
  reg [31:0] _RAND_550;
  reg [31:0] _RAND_551;
  reg [31:0] _RAND_552;
  reg [31:0] _RAND_553;
  reg [31:0] _RAND_554;
  reg [31:0] _RAND_555;
  reg [31:0] _RAND_556;
  reg [31:0] _RAND_557;
  reg [31:0] _RAND_558;
  reg [31:0] _RAND_559;
  reg [31:0] _RAND_560;
  reg [31:0] _RAND_561;
  reg [31:0] _RAND_562;
  reg [31:0] _RAND_563;
  reg [31:0] _RAND_564;
  reg [31:0] _RAND_565;
  reg [31:0] _RAND_566;
  reg [31:0] _RAND_567;
  reg [31:0] _RAND_568;
  reg [31:0] _RAND_569;
  reg [31:0] _RAND_570;
  reg [31:0] _RAND_571;
  reg [31:0] _RAND_572;
  reg [31:0] _RAND_573;
  reg [31:0] _RAND_574;
  reg [31:0] _RAND_575;
  reg [31:0] _RAND_576;
  reg [31:0] _RAND_577;
  reg [31:0] _RAND_578;
  reg [31:0] _RAND_579;
  reg [31:0] _RAND_580;
  reg [31:0] _RAND_581;
  reg [31:0] _RAND_582;
  reg [31:0] _RAND_583;
  reg [31:0] _RAND_584;
  reg [31:0] _RAND_585;
  reg [31:0] _RAND_586;
  reg [31:0] _RAND_587;
  reg [31:0] _RAND_588;
  reg [31:0] _RAND_589;
  reg [31:0] _RAND_590;
  reg [31:0] _RAND_591;
  reg [31:0] _RAND_592;
  reg [31:0] _RAND_593;
  reg [31:0] _RAND_594;
  reg [31:0] _RAND_595;
  reg [31:0] _RAND_596;
  reg [31:0] _RAND_597;
  reg [31:0] _RAND_598;
  reg [31:0] _RAND_599;
  reg [31:0] _RAND_600;
  reg [31:0] _RAND_601;
  reg [31:0] _RAND_602;
  reg [31:0] _RAND_603;
  reg [31:0] _RAND_604;
  reg [31:0] _RAND_605;
  reg [31:0] _RAND_606;
  reg [31:0] _RAND_607;
  reg [31:0] _RAND_608;
  reg [31:0] _RAND_609;
  reg [31:0] _RAND_610;
  reg [31:0] _RAND_611;
  reg [31:0] _RAND_612;
  reg [31:0] _RAND_613;
  reg [31:0] _RAND_614;
  reg [31:0] _RAND_615;
  reg [31:0] _RAND_616;
  reg [31:0] _RAND_617;
  reg [31:0] _RAND_618;
  reg [31:0] _RAND_619;
  reg [31:0] _RAND_620;
  reg [31:0] _RAND_621;
  reg [31:0] _RAND_622;
  reg [31:0] _RAND_623;
  reg [31:0] _RAND_624;
  reg [31:0] _RAND_625;
  reg [31:0] _RAND_626;
  reg [31:0] _RAND_627;
  reg [31:0] _RAND_628;
  reg [31:0] _RAND_629;
  reg [31:0] _RAND_630;
  reg [31:0] _RAND_631;
  reg [31:0] _RAND_632;
  reg [31:0] _RAND_633;
  reg [31:0] _RAND_634;
  reg [31:0] _RAND_635;
  reg [31:0] _RAND_636;
  reg [31:0] _RAND_637;
  reg [31:0] _RAND_638;
  reg [31:0] _RAND_639;
  reg [31:0] _RAND_640;
  reg [31:0] _RAND_641;
  reg [31:0] _RAND_642;
  reg [31:0] _RAND_643;
  reg [31:0] _RAND_644;
  reg [31:0] _RAND_645;
  reg [31:0] _RAND_646;
  reg [31:0] _RAND_647;
  reg [31:0] _RAND_648;
  reg [31:0] _RAND_649;
  reg [31:0] _RAND_650;
  reg [31:0] _RAND_651;
  reg [31:0] _RAND_652;
  reg [31:0] _RAND_653;
  reg [31:0] _RAND_654;
  reg [31:0] _RAND_655;
  reg [31:0] _RAND_656;
  reg [31:0] _RAND_657;
  reg [31:0] _RAND_658;
  reg [31:0] _RAND_659;
  reg [31:0] _RAND_660;
  reg [31:0] _RAND_661;
  reg [31:0] _RAND_662;
  reg [31:0] _RAND_663;
  reg [31:0] _RAND_664;
  reg [31:0] _RAND_665;
  reg [31:0] _RAND_666;
  reg [31:0] _RAND_667;
  reg [31:0] _RAND_668;
  reg [31:0] _RAND_669;
  reg [31:0] _RAND_670;
  reg [31:0] _RAND_671;
  reg [31:0] _RAND_672;
  reg [31:0] _RAND_673;
  reg [31:0] _RAND_674;
  reg [31:0] _RAND_675;
  reg [31:0] _RAND_676;
  reg [31:0] _RAND_677;
  reg [31:0] _RAND_678;
  reg [31:0] _RAND_679;
  reg [31:0] _RAND_680;
  reg [31:0] _RAND_681;
  reg [31:0] _RAND_682;
  reg [31:0] _RAND_683;
  reg [31:0] _RAND_684;
  reg [31:0] _RAND_685;
  reg [31:0] _RAND_686;
  reg [31:0] _RAND_687;
  reg [31:0] _RAND_688;
  reg [31:0] _RAND_689;
  reg [31:0] _RAND_690;
  reg [31:0] _RAND_691;
  reg [31:0] _RAND_692;
  reg [31:0] _RAND_693;
  reg [31:0] _RAND_694;
  reg [31:0] _RAND_695;
  reg [31:0] _RAND_696;
  reg [31:0] _RAND_697;
  reg [31:0] _RAND_698;
  reg [31:0] _RAND_699;
  reg [31:0] _RAND_700;
  reg [31:0] _RAND_701;
  reg [31:0] _RAND_702;
  reg [31:0] _RAND_703;
  reg [31:0] _RAND_704;
  reg [31:0] _RAND_705;
  reg [31:0] _RAND_706;
  reg [31:0] _RAND_707;
  reg [31:0] _RAND_708;
  reg [31:0] _RAND_709;
  reg [31:0] _RAND_710;
  reg [31:0] _RAND_711;
  reg [31:0] _RAND_712;
  reg [31:0] _RAND_713;
  reg [31:0] _RAND_714;
  reg [31:0] _RAND_715;
  reg [31:0] _RAND_716;
  reg [31:0] _RAND_717;
  reg [31:0] _RAND_718;
  reg [31:0] _RAND_719;
  reg [31:0] _RAND_720;
  reg [31:0] _RAND_721;
  reg [31:0] _RAND_722;
  reg [31:0] _RAND_723;
  reg [31:0] _RAND_724;
  reg [31:0] _RAND_725;
  reg [31:0] _RAND_726;
  reg [31:0] _RAND_727;
  reg [31:0] _RAND_728;
  reg [31:0] _RAND_729;
  reg [31:0] _RAND_730;
  reg [31:0] _RAND_731;
  reg [31:0] _RAND_732;
  reg [31:0] _RAND_733;
  reg [31:0] _RAND_734;
  reg [31:0] _RAND_735;
  reg [31:0] _RAND_736;
  reg [31:0] _RAND_737;
  reg [31:0] _RAND_738;
  reg [31:0] _RAND_739;
  reg [31:0] _RAND_740;
  reg [31:0] _RAND_741;
  reg [31:0] _RAND_742;
  reg [31:0] _RAND_743;
  reg [31:0] _RAND_744;
  reg [31:0] _RAND_745;
  reg [31:0] _RAND_746;
  reg [31:0] _RAND_747;
  reg [31:0] _RAND_748;
  reg [31:0] _RAND_749;
  reg [31:0] _RAND_750;
  reg [31:0] _RAND_751;
  reg [31:0] _RAND_752;
  reg [31:0] _RAND_753;
  reg [31:0] _RAND_754;
  reg [31:0] _RAND_755;
  reg [31:0] _RAND_756;
  reg [31:0] _RAND_757;
  reg [31:0] _RAND_758;
  reg [31:0] _RAND_759;
  reg [31:0] _RAND_760;
  reg [31:0] _RAND_761;
  reg [31:0] _RAND_762;
  reg [31:0] _RAND_763;
  reg [31:0] _RAND_764;
  reg [31:0] _RAND_765;
  reg [31:0] _RAND_766;
  reg [31:0] _RAND_767;
  reg [31:0] _RAND_768;
  reg [31:0] _RAND_769;
  reg [31:0] _RAND_770;
  reg [31:0] _RAND_771;
  reg [31:0] _RAND_772;
  reg [31:0] _RAND_773;
  reg [31:0] _RAND_774;
  reg [31:0] _RAND_775;
  reg [31:0] _RAND_776;
  reg [31:0] _RAND_777;
  reg [31:0] _RAND_778;
  reg [31:0] _RAND_779;
  reg [31:0] _RAND_780;
  reg [31:0] _RAND_781;
  reg [31:0] _RAND_782;
  reg [31:0] _RAND_783;
`endif // RANDOMIZE_REG_INIT
  wire [15:0] SMulAdd_io_a_1; // @[ChiselImProc.scala 300:30]
  wire [15:0] SMulAdd_io_a_2; // @[ChiselImProc.scala 300:30]
  wire [15:0] SMulAdd_io_a_3; // @[ChiselImProc.scala 300:30]
  wire [15:0] SMulAdd_io_a_5; // @[ChiselImProc.scala 300:30]
  wire [15:0] SMulAdd_io_a_6; // @[ChiselImProc.scala 300:30]
  wire [15:0] SMulAdd_io_a_7; // @[ChiselImProc.scala 300:30]
  wire [15:0] SMulAdd_io_b_0; // @[ChiselImProc.scala 300:30]
  wire [15:0] SMulAdd_io_b_1; // @[ChiselImProc.scala 300:30]
  wire [15:0] SMulAdd_io_b_2; // @[ChiselImProc.scala 300:30]
  wire [15:0] SMulAdd_io_b_3; // @[ChiselImProc.scala 300:30]
  wire [15:0] SMulAdd_io_b_4; // @[ChiselImProc.scala 300:30]
  wire [15:0] SMulAdd_io_b_5; // @[ChiselImProc.scala 300:30]
  wire [15:0] SMulAdd_io_b_6; // @[ChiselImProc.scala 300:30]
  wire [15:0] SMulAdd_io_b_7; // @[ChiselImProc.scala 300:30]
  wire [15:0] SMulAdd_io_b_8; // @[ChiselImProc.scala 300:30]
  wire [31:0] SMulAdd_io_output; // @[ChiselImProc.scala 300:30]
  wire [15:0] SMulAdd_1_io_a_1; // @[ChiselImProc.scala 301:30]
  wire [15:0] SMulAdd_1_io_a_2; // @[ChiselImProc.scala 301:30]
  wire [15:0] SMulAdd_1_io_a_3; // @[ChiselImProc.scala 301:30]
  wire [15:0] SMulAdd_1_io_a_5; // @[ChiselImProc.scala 301:30]
  wire [15:0] SMulAdd_1_io_a_6; // @[ChiselImProc.scala 301:30]
  wire [15:0] SMulAdd_1_io_a_7; // @[ChiselImProc.scala 301:30]
  wire [15:0] SMulAdd_1_io_b_0; // @[ChiselImProc.scala 301:30]
  wire [15:0] SMulAdd_1_io_b_1; // @[ChiselImProc.scala 301:30]
  wire [15:0] SMulAdd_1_io_b_2; // @[ChiselImProc.scala 301:30]
  wire [15:0] SMulAdd_1_io_b_3; // @[ChiselImProc.scala 301:30]
  wire [15:0] SMulAdd_1_io_b_4; // @[ChiselImProc.scala 301:30]
  wire [15:0] SMulAdd_1_io_b_5; // @[ChiselImProc.scala 301:30]
  wire [15:0] SMulAdd_1_io_b_6; // @[ChiselImProc.scala 301:30]
  wire [15:0] SMulAdd_1_io_b_7; // @[ChiselImProc.scala 301:30]
  wire [15:0] SMulAdd_1_io_b_8; // @[ChiselImProc.scala 301:30]
  wire [31:0] SMulAdd_1_io_output; // @[ChiselImProc.scala 301:30]
  wire [31:0] SqrtExtractionUInt_io_z; // @[ChiselImProc.scala 314:35]
  wire [15:0] SqrtExtractionUInt_io_q; // @[ChiselImProc.scala 314:35]
  reg [1:0] stateReg; // @[ChiselImProc.scala 62:28]
  reg [7:0] dataReg; // @[ChiselImProc.scala 64:23]
  reg [7:0] shadowReg; // @[ChiselImProc.scala 66:25]
  reg  userReg; // @[ChiselImProc.scala 67:23]
  reg  shadowUserReg; // @[ChiselImProc.scala 68:29]
  reg  lastReg; // @[ChiselImProc.scala 69:23]
  reg  shadowLastReg; // @[ChiselImProc.scala 70:29]
  reg [7:0] lineBuffer_0; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_1; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_2; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_3; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_4; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_5; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_6; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_7; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_8; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_9; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_10; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_11; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_12; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_13; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_14; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_15; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_16; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_17; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_18; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_19; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_20; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_21; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_22; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_23; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_24; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_25; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_26; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_27; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_28; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_29; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_30; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_31; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_32; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_33; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_34; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_35; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_36; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_37; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_38; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_39; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_40; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_41; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_42; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_43; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_44; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_45; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_46; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_47; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_48; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_49; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_50; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_51; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_52; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_53; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_54; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_55; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_56; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_57; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_58; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_59; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_60; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_61; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_62; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_63; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_64; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_65; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_66; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_67; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_68; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_69; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_70; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_71; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_72; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_73; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_74; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_75; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_76; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_77; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_78; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_79; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_80; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_81; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_82; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_83; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_84; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_85; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_86; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_87; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_88; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_89; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_90; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_91; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_92; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_93; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_94; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_95; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_96; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_97; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_98; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_99; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_100; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_101; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_102; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_103; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_104; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_105; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_106; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_107; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_108; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_109; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_110; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_111; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_112; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_113; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_114; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_115; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_116; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_117; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_118; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_119; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_120; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_121; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_122; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_123; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_124; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_125; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_126; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_127; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_128; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_129; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_130; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_131; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_132; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_133; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_134; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_135; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_136; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_137; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_138; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_139; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_140; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_141; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_142; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_143; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_144; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_145; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_146; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_147; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_148; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_149; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_150; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_151; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_152; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_153; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_154; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_155; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_156; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_157; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_158; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_159; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_160; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_161; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_162; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_163; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_164; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_165; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_166; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_167; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_168; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_169; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_170; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_171; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_172; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_173; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_174; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_175; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_176; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_177; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_178; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_179; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_180; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_181; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_182; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_183; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_184; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_185; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_186; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_187; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_188; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_189; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_190; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_191; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_192; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_193; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_194; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_195; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_196; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_197; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_198; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_199; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_200; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_201; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_202; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_203; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_204; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_205; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_206; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_207; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_208; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_209; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_210; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_211; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_212; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_213; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_214; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_215; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_216; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_217; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_218; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_219; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_220; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_221; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_222; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_223; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_224; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_225; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_226; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_227; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_228; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_229; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_230; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_231; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_232; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_233; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_234; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_235; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_236; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_237; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_238; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_239; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_240; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_241; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_242; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_243; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_244; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_245; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_246; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_247; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_248; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_249; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_250; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_251; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_252; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_253; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_254; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_255; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_256; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_257; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_258; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_259; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_260; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_261; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_262; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_263; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_264; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_265; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_266; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_267; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_268; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_269; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_270; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_271; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_272; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_273; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_274; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_275; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_276; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_277; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_278; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_279; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_280; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_281; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_282; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_283; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_284; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_285; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_286; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_287; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_288; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_289; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_290; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_291; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_292; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_293; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_294; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_295; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_296; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_297; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_298; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_299; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_300; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_301; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_302; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_303; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_304; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_305; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_306; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_307; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_308; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_309; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_310; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_311; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_312; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_313; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_314; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_315; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_316; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_317; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_318; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_319; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_320; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_321; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_322; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_323; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_324; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_325; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_326; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_327; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_328; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_329; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_330; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_331; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_332; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_333; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_334; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_335; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_336; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_337; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_338; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_339; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_340; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_341; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_342; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_343; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_344; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_345; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_346; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_347; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_348; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_349; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_350; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_351; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_352; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_353; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_354; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_355; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_356; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_357; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_358; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_359; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_360; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_361; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_362; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_363; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_364; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_365; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_366; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_367; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_368; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_369; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_370; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_371; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_372; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_373; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_374; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_375; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_376; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_377; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_378; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_379; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_380; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_381; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_382; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_383; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_384; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_385; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_386; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_387; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_388; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_389; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_390; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_391; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_392; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_393; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_394; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_395; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_396; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_397; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_398; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_399; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_400; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_401; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_402; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_403; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_404; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_405; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_406; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_407; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_408; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_409; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_410; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_411; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_412; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_413; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_414; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_415; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_416; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_417; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_418; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_419; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_420; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_421; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_422; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_423; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_424; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_425; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_426; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_427; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_428; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_429; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_430; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_431; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_432; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_433; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_434; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_435; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_436; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_437; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_438; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_439; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_440; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_441; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_442; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_443; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_444; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_445; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_446; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_447; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_448; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_449; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_450; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_451; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_452; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_453; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_454; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_455; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_456; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_457; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_458; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_459; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_460; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_461; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_462; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_463; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_464; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_465; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_466; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_467; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_468; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_469; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_470; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_471; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_472; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_473; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_474; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_475; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_476; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_477; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_478; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_479; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_480; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_481; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_482; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_483; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_484; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_485; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_486; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_487; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_488; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_489; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_490; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_491; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_492; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_493; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_494; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_495; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_496; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_497; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_498; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_499; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_500; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_501; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_502; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_503; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_504; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_505; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_506; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_507; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_508; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_509; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_510; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_511; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_512; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_513; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_514; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_515; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_516; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_517; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_518; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_519; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_520; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_521; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_522; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_523; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_524; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_525; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_526; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_527; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_528; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_529; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_530; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_531; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_532; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_533; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_534; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_535; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_536; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_537; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_538; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_539; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_540; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_541; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_542; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_543; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_544; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_545; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_546; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_547; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_548; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_549; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_550; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_551; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_552; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_553; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_554; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_555; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_556; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_557; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_558; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_559; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_560; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_561; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_562; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_563; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_564; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_565; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_566; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_567; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_568; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_569; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_570; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_571; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_572; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_573; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_574; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_575; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_576; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_577; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_578; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_579; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_580; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_581; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_582; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_583; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_584; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_585; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_586; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_587; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_588; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_589; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_590; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_591; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_592; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_593; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_594; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_595; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_596; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_597; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_598; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_599; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_600; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_601; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_602; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_603; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_604; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_605; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_606; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_607; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_608; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_609; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_610; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_611; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_612; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_613; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_614; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_615; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_616; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_617; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_618; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_619; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_620; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_621; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_622; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_623; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_624; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_625; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_626; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_627; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_628; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_629; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_630; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_631; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_632; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_633; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_634; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_635; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_636; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_637; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_638; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_639; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_640; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_641; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_642; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_643; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_644; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_645; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_646; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_647; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_648; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_649; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_650; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_651; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_652; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_653; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_654; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_655; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_656; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_657; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_658; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_659; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_660; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_661; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_662; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_663; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_664; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_665; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_666; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_667; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_668; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_669; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_670; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_671; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_672; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_673; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_674; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_675; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_676; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_677; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_678; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_679; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_680; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_681; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_682; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_683; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_684; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_685; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_686; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_687; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_688; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_689; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_690; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_691; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_692; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_693; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_694; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_695; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_696; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_697; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_698; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_699; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_700; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_701; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_702; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_703; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_704; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_705; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_706; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_707; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_708; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_709; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_710; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_711; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_712; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_713; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_714; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_715; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_716; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_717; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_718; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_719; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_720; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_721; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_722; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_723; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_724; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_725; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_726; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_727; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_728; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_729; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_730; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_731; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_732; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_733; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_734; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_735; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_736; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_737; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_738; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_739; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_740; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_741; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_742; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_743; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_744; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_745; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_746; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_747; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_748; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_749; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_750; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_751; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_752; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_753; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_754; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_755; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_756; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_757; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_758; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_759; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_760; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_761; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_762; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_763; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_764; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_765; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_766; // @[ChiselImProc.scala 280:26]
  reg [7:0] lineBuffer_767; // @[ChiselImProc.scala 280:26]
  reg [15:0] windowBuffer_0; // @[ChiselImProc.scala 281:28]
  reg [15:0] windowBuffer_1; // @[ChiselImProc.scala 281:28]
  reg [15:0] windowBuffer_2; // @[ChiselImProc.scala 281:28]
  reg [15:0] windowBuffer_3; // @[ChiselImProc.scala 281:28]
  reg [15:0] windowBuffer_4; // @[ChiselImProc.scala 281:28]
  reg [15:0] windowBuffer_5; // @[ChiselImProc.scala 281:28]
  reg [15:0] windowBuffer_6; // @[ChiselImProc.scala 281:28]
  reg [15:0] windowBuffer_7; // @[ChiselImProc.scala 281:28]
  reg [15:0] windowBuffer_8; // @[ChiselImProc.scala 281:28]
  wire  _T = 2'h0 == stateReg; // @[Conditional.scala 37:30]
  wire  _T_1 = 2'h1 == stateReg; // @[Conditional.scala 37:30]
  wire  _T_2 = ~io_enq_valid; // @[ChiselImProc.scala 84:39]
  wire  _T_3 = io_deq_ready & _T_2; // @[ChiselImProc.scala 84:36]
  wire  _T_4 = io_deq_ready & io_enq_valid; // @[ChiselImProc.scala 87:42]
  wire  _T_5 = ~io_deq_ready; // @[ChiselImProc.scala 92:29]
  wire  _T_6 = _T_5 & io_enq_valid; // @[ChiselImProc.scala 92:43]
  wire  _T_7 = 2'h2 == stateReg; // @[Conditional.scala 37:30]
  wire  _T_8 = 2'h3 == stateReg; // @[Conditional.scala 37:30]
  wire  _T_9 = stateReg == 2'h0; // @[ChiselImProc.scala 116:35]
  wire  _T_10 = stateReg == 2'h1; // @[ChiselImProc.scala 116:57]
  wire  _T_11 = _T_9 | _T_10; // @[ChiselImProc.scala 116:45]
  wire  _T_12 = stateReg == 2'h3; // @[ChiselImProc.scala 116:77]
  wire  _T_15 = stateReg == 2'h2; // @[ChiselImProc.scala 117:55]
  wire  _T_16 = _T_10 | _T_15; // @[ChiselImProc.scala 117:43]
  wire  sel = _T_16 & io_deq_ready; // @[ChiselImProc.scala 286:47]
  wire [16:0] _T_795 = {{9'd0}, lineBuffer_255}; // @[ChiselImProc.scala 297:80]
  wire [15:0] _T_797 = _T_795[15:0]; // @[ChiselImProc.scala 297:110]
  wire [16:0] _T_799 = {{9'd0}, lineBuffer_511}; // @[ChiselImProc.scala 297:80]
  wire [15:0] _T_801 = _T_799[15:0]; // @[ChiselImProc.scala 297:110]
  wire [16:0] _T_803 = {{9'd0}, lineBuffer_767}; // @[ChiselImProc.scala 297:80]
  wire [15:0] _T_805 = _T_803[15:0]; // @[ChiselImProc.scala 297:110]
  wire [63:0] _T_807 = $signed(SMulAdd_io_output) * $signed(SMulAdd_io_output); // @[ChiselImProc.scala 311:30]
  wire [63:0] _T_808 = $signed(SMulAdd_1_io_output) * $signed(SMulAdd_1_io_output); // @[ChiselImProc.scala 311:60]
  wire [63:0] _T_812 = $signed(_T_807) + $signed(_T_808); // @[ChiselImProc.scala 311:76]
  wire [15:0] pix_sqrt_euc = SqrtExtractionUInt_io_q; // @[ChiselImProc.scala 309:28 ChiselImProc.scala 316:18]
  wire  _T_813 = pix_sqrt_euc > 16'hff; // @[ChiselImProc.scala 318:36]
  wire [15:0] pix_sobel = _T_813 ? 16'hff : pix_sqrt_euc; // @[ChiselImProc.scala 318:22]
  wire  _T_815 = $signed(SMulAdd_io_output) == 32'sh0; // @[ChiselImProc.scala 321:33]
  wire [41:0] _T_816 = $signed(SMulAdd_1_io_output) * 32'sh100; // @[ChiselImProc.scala 321:70]
  wire [41:0] _GEN_47 = {{10{SMulAdd_io_output[31]}},SMulAdd_io_output}; // @[ChiselImProc.scala 321:80]
  wire [42:0] _T_817 = $signed(_T_816) / $signed(_GEN_47); // @[ChiselImProc.scala 321:80]
  wire [42:0] _T_818 = _T_815 ? $signed(43'sh7fffffff) : $signed(_T_817); // @[ChiselImProc.scala 321:18]
  wire [31:0] t_int = _T_818[31:0]; // @[ChiselImProc.scala 320:22 ChiselImProc.scala 321:11]
  wire  _T_819 = -32'sh26a < $signed(t_int); // @[ChiselImProc.scala 324:18]
  wire  _T_820 = $signed(t_int) <= -32'sh6a; // @[ChiselImProc.scala 324:35]
  wire  _T_821 = _T_819 & _T_820; // @[ChiselImProc.scala 324:26]
  wire  _T_822 = -32'sh6a < $signed(t_int); // @[ChiselImProc.scala 326:24]
  wire  _T_823 = $signed(t_int) <= 32'sh6a; // @[ChiselImProc.scala 326:41]
  wire  _T_824 = _T_822 & _T_823; // @[ChiselImProc.scala 326:32]
  wire  _T_825 = 32'sh6a < $signed(t_int); // @[ChiselImProc.scala 328:23]
  wire  _T_826 = $signed(t_int) <= 32'sh26a; // @[ChiselImProc.scala 328:40]
  wire  _T_827 = _T_825 & _T_826; // @[ChiselImProc.scala 328:31]
  wire [1:0] _GEN_44 = _T_827 ? 2'h1 : 2'h2; // @[ChiselImProc.scala 328:50]
  wire [1:0] _GEN_45 = _T_824 ? 2'h0 : _GEN_44; // @[ChiselImProc.scala 326:51]
  SMulAdd SMulAdd ( // @[ChiselImProc.scala 300:30]
    .io_a_1(SMulAdd_io_a_1),
    .io_a_2(SMulAdd_io_a_2),
    .io_a_3(SMulAdd_io_a_3),
    .io_a_5(SMulAdd_io_a_5),
    .io_a_6(SMulAdd_io_a_6),
    .io_a_7(SMulAdd_io_a_7),
    .io_b_0(SMulAdd_io_b_0),
    .io_b_1(SMulAdd_io_b_1),
    .io_b_2(SMulAdd_io_b_2),
    .io_b_3(SMulAdd_io_b_3),
    .io_b_4(SMulAdd_io_b_4),
    .io_b_5(SMulAdd_io_b_5),
    .io_b_6(SMulAdd_io_b_6),
    .io_b_7(SMulAdd_io_b_7),
    .io_b_8(SMulAdd_io_b_8),
    .io_output(SMulAdd_io_output)
  );
  SMulAdd SMulAdd_1 ( // @[ChiselImProc.scala 301:30]
    .io_a_1(SMulAdd_1_io_a_1),
    .io_a_2(SMulAdd_1_io_a_2),
    .io_a_3(SMulAdd_1_io_a_3),
    .io_a_5(SMulAdd_1_io_a_5),
    .io_a_6(SMulAdd_1_io_a_6),
    .io_a_7(SMulAdd_1_io_a_7),
    .io_b_0(SMulAdd_1_io_b_0),
    .io_b_1(SMulAdd_1_io_b_1),
    .io_b_2(SMulAdd_1_io_b_2),
    .io_b_3(SMulAdd_1_io_b_3),
    .io_b_4(SMulAdd_1_io_b_4),
    .io_b_5(SMulAdd_1_io_b_5),
    .io_b_6(SMulAdd_1_io_b_6),
    .io_b_7(SMulAdd_1_io_b_7),
    .io_b_8(SMulAdd_1_io_b_8),
    .io_output(SMulAdd_1_io_output)
  );
  SqrtExtractionUInt SqrtExtractionUInt ( // @[ChiselImProc.scala 314:35]
    .io_z(SqrtExtractionUInt_io_z),
    .io_q(SqrtExtractionUInt_io_q)
  );
  assign io_enq_ready = _T_11 | _T_12; // @[ChiselImProc.scala 116:22]
  assign io_deq_valid = _T_10 | _T_15; // @[ChiselImProc.scala 117:22]
  assign io_deq_bits_grad_dir = _T_821 ? 2'h3 : _GEN_45; // @[ChiselImProc.scala 334:26]
  assign io_deq_bits_value = pix_sobel[7:0]; // @[ChiselImProc.scala 335:23]
  assign io_deq_user = userReg; // @[ChiselImProc.scala 114:21]
  assign io_deq_last = lastReg; // @[ChiselImProc.scala 113:21]
  assign SMulAdd_io_a_1 = 16'sh0; // @[ChiselImProc.scala 303:14]
  assign SMulAdd_io_a_2 = -16'sh1; // @[ChiselImProc.scala 303:14]
  assign SMulAdd_io_a_3 = 16'sh2; // @[ChiselImProc.scala 303:14]
  assign SMulAdd_io_a_5 = -16'sh2; // @[ChiselImProc.scala 303:14]
  assign SMulAdd_io_a_6 = 16'sh1; // @[ChiselImProc.scala 303:14]
  assign SMulAdd_io_a_7 = 16'sh0; // @[ChiselImProc.scala 303:14]
  assign SMulAdd_io_b_0 = windowBuffer_0; // @[ChiselImProc.scala 304:14]
  assign SMulAdd_io_b_1 = windowBuffer_1; // @[ChiselImProc.scala 304:14]
  assign SMulAdd_io_b_2 = windowBuffer_2; // @[ChiselImProc.scala 304:14]
  assign SMulAdd_io_b_3 = windowBuffer_3; // @[ChiselImProc.scala 304:14]
  assign SMulAdd_io_b_4 = windowBuffer_4; // @[ChiselImProc.scala 304:14]
  assign SMulAdd_io_b_5 = windowBuffer_5; // @[ChiselImProc.scala 304:14]
  assign SMulAdd_io_b_6 = windowBuffer_6; // @[ChiselImProc.scala 304:14]
  assign SMulAdd_io_b_7 = windowBuffer_7; // @[ChiselImProc.scala 304:14]
  assign SMulAdd_io_b_8 = windowBuffer_8; // @[ChiselImProc.scala 304:14]
  assign SMulAdd_1_io_a_1 = 16'sh2; // @[ChiselImProc.scala 305:14]
  assign SMulAdd_1_io_a_2 = 16'sh1; // @[ChiselImProc.scala 305:14]
  assign SMulAdd_1_io_a_3 = 16'sh0; // @[ChiselImProc.scala 305:14]
  assign SMulAdd_1_io_a_5 = 16'sh0; // @[ChiselImProc.scala 305:14]
  assign SMulAdd_1_io_a_6 = -16'sh1; // @[ChiselImProc.scala 305:14]
  assign SMulAdd_1_io_a_7 = -16'sh2; // @[ChiselImProc.scala 305:14]
  assign SMulAdd_1_io_b_0 = windowBuffer_0; // @[ChiselImProc.scala 306:14]
  assign SMulAdd_1_io_b_1 = windowBuffer_1; // @[ChiselImProc.scala 306:14]
  assign SMulAdd_1_io_b_2 = windowBuffer_2; // @[ChiselImProc.scala 306:14]
  assign SMulAdd_1_io_b_3 = windowBuffer_3; // @[ChiselImProc.scala 306:14]
  assign SMulAdd_1_io_b_4 = windowBuffer_4; // @[ChiselImProc.scala 306:14]
  assign SMulAdd_1_io_b_5 = windowBuffer_5; // @[ChiselImProc.scala 306:14]
  assign SMulAdd_1_io_b_6 = windowBuffer_6; // @[ChiselImProc.scala 306:14]
  assign SMulAdd_1_io_b_7 = windowBuffer_7; // @[ChiselImProc.scala 306:14]
  assign SMulAdd_1_io_b_8 = windowBuffer_8; // @[ChiselImProc.scala 306:14]
  assign SqrtExtractionUInt_io_z = _T_812[31:0]; // @[ChiselImProc.scala 315:19]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  stateReg = _RAND_0[1:0];
  _RAND_1 = {1{`RANDOM}};
  dataReg = _RAND_1[7:0];
  _RAND_2 = {1{`RANDOM}};
  shadowReg = _RAND_2[7:0];
  _RAND_3 = {1{`RANDOM}};
  userReg = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  shadowUserReg = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  lastReg = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  shadowLastReg = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  lineBuffer_0 = _RAND_7[7:0];
  _RAND_8 = {1{`RANDOM}};
  lineBuffer_1 = _RAND_8[7:0];
  _RAND_9 = {1{`RANDOM}};
  lineBuffer_2 = _RAND_9[7:0];
  _RAND_10 = {1{`RANDOM}};
  lineBuffer_3 = _RAND_10[7:0];
  _RAND_11 = {1{`RANDOM}};
  lineBuffer_4 = _RAND_11[7:0];
  _RAND_12 = {1{`RANDOM}};
  lineBuffer_5 = _RAND_12[7:0];
  _RAND_13 = {1{`RANDOM}};
  lineBuffer_6 = _RAND_13[7:0];
  _RAND_14 = {1{`RANDOM}};
  lineBuffer_7 = _RAND_14[7:0];
  _RAND_15 = {1{`RANDOM}};
  lineBuffer_8 = _RAND_15[7:0];
  _RAND_16 = {1{`RANDOM}};
  lineBuffer_9 = _RAND_16[7:0];
  _RAND_17 = {1{`RANDOM}};
  lineBuffer_10 = _RAND_17[7:0];
  _RAND_18 = {1{`RANDOM}};
  lineBuffer_11 = _RAND_18[7:0];
  _RAND_19 = {1{`RANDOM}};
  lineBuffer_12 = _RAND_19[7:0];
  _RAND_20 = {1{`RANDOM}};
  lineBuffer_13 = _RAND_20[7:0];
  _RAND_21 = {1{`RANDOM}};
  lineBuffer_14 = _RAND_21[7:0];
  _RAND_22 = {1{`RANDOM}};
  lineBuffer_15 = _RAND_22[7:0];
  _RAND_23 = {1{`RANDOM}};
  lineBuffer_16 = _RAND_23[7:0];
  _RAND_24 = {1{`RANDOM}};
  lineBuffer_17 = _RAND_24[7:0];
  _RAND_25 = {1{`RANDOM}};
  lineBuffer_18 = _RAND_25[7:0];
  _RAND_26 = {1{`RANDOM}};
  lineBuffer_19 = _RAND_26[7:0];
  _RAND_27 = {1{`RANDOM}};
  lineBuffer_20 = _RAND_27[7:0];
  _RAND_28 = {1{`RANDOM}};
  lineBuffer_21 = _RAND_28[7:0];
  _RAND_29 = {1{`RANDOM}};
  lineBuffer_22 = _RAND_29[7:0];
  _RAND_30 = {1{`RANDOM}};
  lineBuffer_23 = _RAND_30[7:0];
  _RAND_31 = {1{`RANDOM}};
  lineBuffer_24 = _RAND_31[7:0];
  _RAND_32 = {1{`RANDOM}};
  lineBuffer_25 = _RAND_32[7:0];
  _RAND_33 = {1{`RANDOM}};
  lineBuffer_26 = _RAND_33[7:0];
  _RAND_34 = {1{`RANDOM}};
  lineBuffer_27 = _RAND_34[7:0];
  _RAND_35 = {1{`RANDOM}};
  lineBuffer_28 = _RAND_35[7:0];
  _RAND_36 = {1{`RANDOM}};
  lineBuffer_29 = _RAND_36[7:0];
  _RAND_37 = {1{`RANDOM}};
  lineBuffer_30 = _RAND_37[7:0];
  _RAND_38 = {1{`RANDOM}};
  lineBuffer_31 = _RAND_38[7:0];
  _RAND_39 = {1{`RANDOM}};
  lineBuffer_32 = _RAND_39[7:0];
  _RAND_40 = {1{`RANDOM}};
  lineBuffer_33 = _RAND_40[7:0];
  _RAND_41 = {1{`RANDOM}};
  lineBuffer_34 = _RAND_41[7:0];
  _RAND_42 = {1{`RANDOM}};
  lineBuffer_35 = _RAND_42[7:0];
  _RAND_43 = {1{`RANDOM}};
  lineBuffer_36 = _RAND_43[7:0];
  _RAND_44 = {1{`RANDOM}};
  lineBuffer_37 = _RAND_44[7:0];
  _RAND_45 = {1{`RANDOM}};
  lineBuffer_38 = _RAND_45[7:0];
  _RAND_46 = {1{`RANDOM}};
  lineBuffer_39 = _RAND_46[7:0];
  _RAND_47 = {1{`RANDOM}};
  lineBuffer_40 = _RAND_47[7:0];
  _RAND_48 = {1{`RANDOM}};
  lineBuffer_41 = _RAND_48[7:0];
  _RAND_49 = {1{`RANDOM}};
  lineBuffer_42 = _RAND_49[7:0];
  _RAND_50 = {1{`RANDOM}};
  lineBuffer_43 = _RAND_50[7:0];
  _RAND_51 = {1{`RANDOM}};
  lineBuffer_44 = _RAND_51[7:0];
  _RAND_52 = {1{`RANDOM}};
  lineBuffer_45 = _RAND_52[7:0];
  _RAND_53 = {1{`RANDOM}};
  lineBuffer_46 = _RAND_53[7:0];
  _RAND_54 = {1{`RANDOM}};
  lineBuffer_47 = _RAND_54[7:0];
  _RAND_55 = {1{`RANDOM}};
  lineBuffer_48 = _RAND_55[7:0];
  _RAND_56 = {1{`RANDOM}};
  lineBuffer_49 = _RAND_56[7:0];
  _RAND_57 = {1{`RANDOM}};
  lineBuffer_50 = _RAND_57[7:0];
  _RAND_58 = {1{`RANDOM}};
  lineBuffer_51 = _RAND_58[7:0];
  _RAND_59 = {1{`RANDOM}};
  lineBuffer_52 = _RAND_59[7:0];
  _RAND_60 = {1{`RANDOM}};
  lineBuffer_53 = _RAND_60[7:0];
  _RAND_61 = {1{`RANDOM}};
  lineBuffer_54 = _RAND_61[7:0];
  _RAND_62 = {1{`RANDOM}};
  lineBuffer_55 = _RAND_62[7:0];
  _RAND_63 = {1{`RANDOM}};
  lineBuffer_56 = _RAND_63[7:0];
  _RAND_64 = {1{`RANDOM}};
  lineBuffer_57 = _RAND_64[7:0];
  _RAND_65 = {1{`RANDOM}};
  lineBuffer_58 = _RAND_65[7:0];
  _RAND_66 = {1{`RANDOM}};
  lineBuffer_59 = _RAND_66[7:0];
  _RAND_67 = {1{`RANDOM}};
  lineBuffer_60 = _RAND_67[7:0];
  _RAND_68 = {1{`RANDOM}};
  lineBuffer_61 = _RAND_68[7:0];
  _RAND_69 = {1{`RANDOM}};
  lineBuffer_62 = _RAND_69[7:0];
  _RAND_70 = {1{`RANDOM}};
  lineBuffer_63 = _RAND_70[7:0];
  _RAND_71 = {1{`RANDOM}};
  lineBuffer_64 = _RAND_71[7:0];
  _RAND_72 = {1{`RANDOM}};
  lineBuffer_65 = _RAND_72[7:0];
  _RAND_73 = {1{`RANDOM}};
  lineBuffer_66 = _RAND_73[7:0];
  _RAND_74 = {1{`RANDOM}};
  lineBuffer_67 = _RAND_74[7:0];
  _RAND_75 = {1{`RANDOM}};
  lineBuffer_68 = _RAND_75[7:0];
  _RAND_76 = {1{`RANDOM}};
  lineBuffer_69 = _RAND_76[7:0];
  _RAND_77 = {1{`RANDOM}};
  lineBuffer_70 = _RAND_77[7:0];
  _RAND_78 = {1{`RANDOM}};
  lineBuffer_71 = _RAND_78[7:0];
  _RAND_79 = {1{`RANDOM}};
  lineBuffer_72 = _RAND_79[7:0];
  _RAND_80 = {1{`RANDOM}};
  lineBuffer_73 = _RAND_80[7:0];
  _RAND_81 = {1{`RANDOM}};
  lineBuffer_74 = _RAND_81[7:0];
  _RAND_82 = {1{`RANDOM}};
  lineBuffer_75 = _RAND_82[7:0];
  _RAND_83 = {1{`RANDOM}};
  lineBuffer_76 = _RAND_83[7:0];
  _RAND_84 = {1{`RANDOM}};
  lineBuffer_77 = _RAND_84[7:0];
  _RAND_85 = {1{`RANDOM}};
  lineBuffer_78 = _RAND_85[7:0];
  _RAND_86 = {1{`RANDOM}};
  lineBuffer_79 = _RAND_86[7:0];
  _RAND_87 = {1{`RANDOM}};
  lineBuffer_80 = _RAND_87[7:0];
  _RAND_88 = {1{`RANDOM}};
  lineBuffer_81 = _RAND_88[7:0];
  _RAND_89 = {1{`RANDOM}};
  lineBuffer_82 = _RAND_89[7:0];
  _RAND_90 = {1{`RANDOM}};
  lineBuffer_83 = _RAND_90[7:0];
  _RAND_91 = {1{`RANDOM}};
  lineBuffer_84 = _RAND_91[7:0];
  _RAND_92 = {1{`RANDOM}};
  lineBuffer_85 = _RAND_92[7:0];
  _RAND_93 = {1{`RANDOM}};
  lineBuffer_86 = _RAND_93[7:0];
  _RAND_94 = {1{`RANDOM}};
  lineBuffer_87 = _RAND_94[7:0];
  _RAND_95 = {1{`RANDOM}};
  lineBuffer_88 = _RAND_95[7:0];
  _RAND_96 = {1{`RANDOM}};
  lineBuffer_89 = _RAND_96[7:0];
  _RAND_97 = {1{`RANDOM}};
  lineBuffer_90 = _RAND_97[7:0];
  _RAND_98 = {1{`RANDOM}};
  lineBuffer_91 = _RAND_98[7:0];
  _RAND_99 = {1{`RANDOM}};
  lineBuffer_92 = _RAND_99[7:0];
  _RAND_100 = {1{`RANDOM}};
  lineBuffer_93 = _RAND_100[7:0];
  _RAND_101 = {1{`RANDOM}};
  lineBuffer_94 = _RAND_101[7:0];
  _RAND_102 = {1{`RANDOM}};
  lineBuffer_95 = _RAND_102[7:0];
  _RAND_103 = {1{`RANDOM}};
  lineBuffer_96 = _RAND_103[7:0];
  _RAND_104 = {1{`RANDOM}};
  lineBuffer_97 = _RAND_104[7:0];
  _RAND_105 = {1{`RANDOM}};
  lineBuffer_98 = _RAND_105[7:0];
  _RAND_106 = {1{`RANDOM}};
  lineBuffer_99 = _RAND_106[7:0];
  _RAND_107 = {1{`RANDOM}};
  lineBuffer_100 = _RAND_107[7:0];
  _RAND_108 = {1{`RANDOM}};
  lineBuffer_101 = _RAND_108[7:0];
  _RAND_109 = {1{`RANDOM}};
  lineBuffer_102 = _RAND_109[7:0];
  _RAND_110 = {1{`RANDOM}};
  lineBuffer_103 = _RAND_110[7:0];
  _RAND_111 = {1{`RANDOM}};
  lineBuffer_104 = _RAND_111[7:0];
  _RAND_112 = {1{`RANDOM}};
  lineBuffer_105 = _RAND_112[7:0];
  _RAND_113 = {1{`RANDOM}};
  lineBuffer_106 = _RAND_113[7:0];
  _RAND_114 = {1{`RANDOM}};
  lineBuffer_107 = _RAND_114[7:0];
  _RAND_115 = {1{`RANDOM}};
  lineBuffer_108 = _RAND_115[7:0];
  _RAND_116 = {1{`RANDOM}};
  lineBuffer_109 = _RAND_116[7:0];
  _RAND_117 = {1{`RANDOM}};
  lineBuffer_110 = _RAND_117[7:0];
  _RAND_118 = {1{`RANDOM}};
  lineBuffer_111 = _RAND_118[7:0];
  _RAND_119 = {1{`RANDOM}};
  lineBuffer_112 = _RAND_119[7:0];
  _RAND_120 = {1{`RANDOM}};
  lineBuffer_113 = _RAND_120[7:0];
  _RAND_121 = {1{`RANDOM}};
  lineBuffer_114 = _RAND_121[7:0];
  _RAND_122 = {1{`RANDOM}};
  lineBuffer_115 = _RAND_122[7:0];
  _RAND_123 = {1{`RANDOM}};
  lineBuffer_116 = _RAND_123[7:0];
  _RAND_124 = {1{`RANDOM}};
  lineBuffer_117 = _RAND_124[7:0];
  _RAND_125 = {1{`RANDOM}};
  lineBuffer_118 = _RAND_125[7:0];
  _RAND_126 = {1{`RANDOM}};
  lineBuffer_119 = _RAND_126[7:0];
  _RAND_127 = {1{`RANDOM}};
  lineBuffer_120 = _RAND_127[7:0];
  _RAND_128 = {1{`RANDOM}};
  lineBuffer_121 = _RAND_128[7:0];
  _RAND_129 = {1{`RANDOM}};
  lineBuffer_122 = _RAND_129[7:0];
  _RAND_130 = {1{`RANDOM}};
  lineBuffer_123 = _RAND_130[7:0];
  _RAND_131 = {1{`RANDOM}};
  lineBuffer_124 = _RAND_131[7:0];
  _RAND_132 = {1{`RANDOM}};
  lineBuffer_125 = _RAND_132[7:0];
  _RAND_133 = {1{`RANDOM}};
  lineBuffer_126 = _RAND_133[7:0];
  _RAND_134 = {1{`RANDOM}};
  lineBuffer_127 = _RAND_134[7:0];
  _RAND_135 = {1{`RANDOM}};
  lineBuffer_128 = _RAND_135[7:0];
  _RAND_136 = {1{`RANDOM}};
  lineBuffer_129 = _RAND_136[7:0];
  _RAND_137 = {1{`RANDOM}};
  lineBuffer_130 = _RAND_137[7:0];
  _RAND_138 = {1{`RANDOM}};
  lineBuffer_131 = _RAND_138[7:0];
  _RAND_139 = {1{`RANDOM}};
  lineBuffer_132 = _RAND_139[7:0];
  _RAND_140 = {1{`RANDOM}};
  lineBuffer_133 = _RAND_140[7:0];
  _RAND_141 = {1{`RANDOM}};
  lineBuffer_134 = _RAND_141[7:0];
  _RAND_142 = {1{`RANDOM}};
  lineBuffer_135 = _RAND_142[7:0];
  _RAND_143 = {1{`RANDOM}};
  lineBuffer_136 = _RAND_143[7:0];
  _RAND_144 = {1{`RANDOM}};
  lineBuffer_137 = _RAND_144[7:0];
  _RAND_145 = {1{`RANDOM}};
  lineBuffer_138 = _RAND_145[7:0];
  _RAND_146 = {1{`RANDOM}};
  lineBuffer_139 = _RAND_146[7:0];
  _RAND_147 = {1{`RANDOM}};
  lineBuffer_140 = _RAND_147[7:0];
  _RAND_148 = {1{`RANDOM}};
  lineBuffer_141 = _RAND_148[7:0];
  _RAND_149 = {1{`RANDOM}};
  lineBuffer_142 = _RAND_149[7:0];
  _RAND_150 = {1{`RANDOM}};
  lineBuffer_143 = _RAND_150[7:0];
  _RAND_151 = {1{`RANDOM}};
  lineBuffer_144 = _RAND_151[7:0];
  _RAND_152 = {1{`RANDOM}};
  lineBuffer_145 = _RAND_152[7:0];
  _RAND_153 = {1{`RANDOM}};
  lineBuffer_146 = _RAND_153[7:0];
  _RAND_154 = {1{`RANDOM}};
  lineBuffer_147 = _RAND_154[7:0];
  _RAND_155 = {1{`RANDOM}};
  lineBuffer_148 = _RAND_155[7:0];
  _RAND_156 = {1{`RANDOM}};
  lineBuffer_149 = _RAND_156[7:0];
  _RAND_157 = {1{`RANDOM}};
  lineBuffer_150 = _RAND_157[7:0];
  _RAND_158 = {1{`RANDOM}};
  lineBuffer_151 = _RAND_158[7:0];
  _RAND_159 = {1{`RANDOM}};
  lineBuffer_152 = _RAND_159[7:0];
  _RAND_160 = {1{`RANDOM}};
  lineBuffer_153 = _RAND_160[7:0];
  _RAND_161 = {1{`RANDOM}};
  lineBuffer_154 = _RAND_161[7:0];
  _RAND_162 = {1{`RANDOM}};
  lineBuffer_155 = _RAND_162[7:0];
  _RAND_163 = {1{`RANDOM}};
  lineBuffer_156 = _RAND_163[7:0];
  _RAND_164 = {1{`RANDOM}};
  lineBuffer_157 = _RAND_164[7:0];
  _RAND_165 = {1{`RANDOM}};
  lineBuffer_158 = _RAND_165[7:0];
  _RAND_166 = {1{`RANDOM}};
  lineBuffer_159 = _RAND_166[7:0];
  _RAND_167 = {1{`RANDOM}};
  lineBuffer_160 = _RAND_167[7:0];
  _RAND_168 = {1{`RANDOM}};
  lineBuffer_161 = _RAND_168[7:0];
  _RAND_169 = {1{`RANDOM}};
  lineBuffer_162 = _RAND_169[7:0];
  _RAND_170 = {1{`RANDOM}};
  lineBuffer_163 = _RAND_170[7:0];
  _RAND_171 = {1{`RANDOM}};
  lineBuffer_164 = _RAND_171[7:0];
  _RAND_172 = {1{`RANDOM}};
  lineBuffer_165 = _RAND_172[7:0];
  _RAND_173 = {1{`RANDOM}};
  lineBuffer_166 = _RAND_173[7:0];
  _RAND_174 = {1{`RANDOM}};
  lineBuffer_167 = _RAND_174[7:0];
  _RAND_175 = {1{`RANDOM}};
  lineBuffer_168 = _RAND_175[7:0];
  _RAND_176 = {1{`RANDOM}};
  lineBuffer_169 = _RAND_176[7:0];
  _RAND_177 = {1{`RANDOM}};
  lineBuffer_170 = _RAND_177[7:0];
  _RAND_178 = {1{`RANDOM}};
  lineBuffer_171 = _RAND_178[7:0];
  _RAND_179 = {1{`RANDOM}};
  lineBuffer_172 = _RAND_179[7:0];
  _RAND_180 = {1{`RANDOM}};
  lineBuffer_173 = _RAND_180[7:0];
  _RAND_181 = {1{`RANDOM}};
  lineBuffer_174 = _RAND_181[7:0];
  _RAND_182 = {1{`RANDOM}};
  lineBuffer_175 = _RAND_182[7:0];
  _RAND_183 = {1{`RANDOM}};
  lineBuffer_176 = _RAND_183[7:0];
  _RAND_184 = {1{`RANDOM}};
  lineBuffer_177 = _RAND_184[7:0];
  _RAND_185 = {1{`RANDOM}};
  lineBuffer_178 = _RAND_185[7:0];
  _RAND_186 = {1{`RANDOM}};
  lineBuffer_179 = _RAND_186[7:0];
  _RAND_187 = {1{`RANDOM}};
  lineBuffer_180 = _RAND_187[7:0];
  _RAND_188 = {1{`RANDOM}};
  lineBuffer_181 = _RAND_188[7:0];
  _RAND_189 = {1{`RANDOM}};
  lineBuffer_182 = _RAND_189[7:0];
  _RAND_190 = {1{`RANDOM}};
  lineBuffer_183 = _RAND_190[7:0];
  _RAND_191 = {1{`RANDOM}};
  lineBuffer_184 = _RAND_191[7:0];
  _RAND_192 = {1{`RANDOM}};
  lineBuffer_185 = _RAND_192[7:0];
  _RAND_193 = {1{`RANDOM}};
  lineBuffer_186 = _RAND_193[7:0];
  _RAND_194 = {1{`RANDOM}};
  lineBuffer_187 = _RAND_194[7:0];
  _RAND_195 = {1{`RANDOM}};
  lineBuffer_188 = _RAND_195[7:0];
  _RAND_196 = {1{`RANDOM}};
  lineBuffer_189 = _RAND_196[7:0];
  _RAND_197 = {1{`RANDOM}};
  lineBuffer_190 = _RAND_197[7:0];
  _RAND_198 = {1{`RANDOM}};
  lineBuffer_191 = _RAND_198[7:0];
  _RAND_199 = {1{`RANDOM}};
  lineBuffer_192 = _RAND_199[7:0];
  _RAND_200 = {1{`RANDOM}};
  lineBuffer_193 = _RAND_200[7:0];
  _RAND_201 = {1{`RANDOM}};
  lineBuffer_194 = _RAND_201[7:0];
  _RAND_202 = {1{`RANDOM}};
  lineBuffer_195 = _RAND_202[7:0];
  _RAND_203 = {1{`RANDOM}};
  lineBuffer_196 = _RAND_203[7:0];
  _RAND_204 = {1{`RANDOM}};
  lineBuffer_197 = _RAND_204[7:0];
  _RAND_205 = {1{`RANDOM}};
  lineBuffer_198 = _RAND_205[7:0];
  _RAND_206 = {1{`RANDOM}};
  lineBuffer_199 = _RAND_206[7:0];
  _RAND_207 = {1{`RANDOM}};
  lineBuffer_200 = _RAND_207[7:0];
  _RAND_208 = {1{`RANDOM}};
  lineBuffer_201 = _RAND_208[7:0];
  _RAND_209 = {1{`RANDOM}};
  lineBuffer_202 = _RAND_209[7:0];
  _RAND_210 = {1{`RANDOM}};
  lineBuffer_203 = _RAND_210[7:0];
  _RAND_211 = {1{`RANDOM}};
  lineBuffer_204 = _RAND_211[7:0];
  _RAND_212 = {1{`RANDOM}};
  lineBuffer_205 = _RAND_212[7:0];
  _RAND_213 = {1{`RANDOM}};
  lineBuffer_206 = _RAND_213[7:0];
  _RAND_214 = {1{`RANDOM}};
  lineBuffer_207 = _RAND_214[7:0];
  _RAND_215 = {1{`RANDOM}};
  lineBuffer_208 = _RAND_215[7:0];
  _RAND_216 = {1{`RANDOM}};
  lineBuffer_209 = _RAND_216[7:0];
  _RAND_217 = {1{`RANDOM}};
  lineBuffer_210 = _RAND_217[7:0];
  _RAND_218 = {1{`RANDOM}};
  lineBuffer_211 = _RAND_218[7:0];
  _RAND_219 = {1{`RANDOM}};
  lineBuffer_212 = _RAND_219[7:0];
  _RAND_220 = {1{`RANDOM}};
  lineBuffer_213 = _RAND_220[7:0];
  _RAND_221 = {1{`RANDOM}};
  lineBuffer_214 = _RAND_221[7:0];
  _RAND_222 = {1{`RANDOM}};
  lineBuffer_215 = _RAND_222[7:0];
  _RAND_223 = {1{`RANDOM}};
  lineBuffer_216 = _RAND_223[7:0];
  _RAND_224 = {1{`RANDOM}};
  lineBuffer_217 = _RAND_224[7:0];
  _RAND_225 = {1{`RANDOM}};
  lineBuffer_218 = _RAND_225[7:0];
  _RAND_226 = {1{`RANDOM}};
  lineBuffer_219 = _RAND_226[7:0];
  _RAND_227 = {1{`RANDOM}};
  lineBuffer_220 = _RAND_227[7:0];
  _RAND_228 = {1{`RANDOM}};
  lineBuffer_221 = _RAND_228[7:0];
  _RAND_229 = {1{`RANDOM}};
  lineBuffer_222 = _RAND_229[7:0];
  _RAND_230 = {1{`RANDOM}};
  lineBuffer_223 = _RAND_230[7:0];
  _RAND_231 = {1{`RANDOM}};
  lineBuffer_224 = _RAND_231[7:0];
  _RAND_232 = {1{`RANDOM}};
  lineBuffer_225 = _RAND_232[7:0];
  _RAND_233 = {1{`RANDOM}};
  lineBuffer_226 = _RAND_233[7:0];
  _RAND_234 = {1{`RANDOM}};
  lineBuffer_227 = _RAND_234[7:0];
  _RAND_235 = {1{`RANDOM}};
  lineBuffer_228 = _RAND_235[7:0];
  _RAND_236 = {1{`RANDOM}};
  lineBuffer_229 = _RAND_236[7:0];
  _RAND_237 = {1{`RANDOM}};
  lineBuffer_230 = _RAND_237[7:0];
  _RAND_238 = {1{`RANDOM}};
  lineBuffer_231 = _RAND_238[7:0];
  _RAND_239 = {1{`RANDOM}};
  lineBuffer_232 = _RAND_239[7:0];
  _RAND_240 = {1{`RANDOM}};
  lineBuffer_233 = _RAND_240[7:0];
  _RAND_241 = {1{`RANDOM}};
  lineBuffer_234 = _RAND_241[7:0];
  _RAND_242 = {1{`RANDOM}};
  lineBuffer_235 = _RAND_242[7:0];
  _RAND_243 = {1{`RANDOM}};
  lineBuffer_236 = _RAND_243[7:0];
  _RAND_244 = {1{`RANDOM}};
  lineBuffer_237 = _RAND_244[7:0];
  _RAND_245 = {1{`RANDOM}};
  lineBuffer_238 = _RAND_245[7:0];
  _RAND_246 = {1{`RANDOM}};
  lineBuffer_239 = _RAND_246[7:0];
  _RAND_247 = {1{`RANDOM}};
  lineBuffer_240 = _RAND_247[7:0];
  _RAND_248 = {1{`RANDOM}};
  lineBuffer_241 = _RAND_248[7:0];
  _RAND_249 = {1{`RANDOM}};
  lineBuffer_242 = _RAND_249[7:0];
  _RAND_250 = {1{`RANDOM}};
  lineBuffer_243 = _RAND_250[7:0];
  _RAND_251 = {1{`RANDOM}};
  lineBuffer_244 = _RAND_251[7:0];
  _RAND_252 = {1{`RANDOM}};
  lineBuffer_245 = _RAND_252[7:0];
  _RAND_253 = {1{`RANDOM}};
  lineBuffer_246 = _RAND_253[7:0];
  _RAND_254 = {1{`RANDOM}};
  lineBuffer_247 = _RAND_254[7:0];
  _RAND_255 = {1{`RANDOM}};
  lineBuffer_248 = _RAND_255[7:0];
  _RAND_256 = {1{`RANDOM}};
  lineBuffer_249 = _RAND_256[7:0];
  _RAND_257 = {1{`RANDOM}};
  lineBuffer_250 = _RAND_257[7:0];
  _RAND_258 = {1{`RANDOM}};
  lineBuffer_251 = _RAND_258[7:0];
  _RAND_259 = {1{`RANDOM}};
  lineBuffer_252 = _RAND_259[7:0];
  _RAND_260 = {1{`RANDOM}};
  lineBuffer_253 = _RAND_260[7:0];
  _RAND_261 = {1{`RANDOM}};
  lineBuffer_254 = _RAND_261[7:0];
  _RAND_262 = {1{`RANDOM}};
  lineBuffer_255 = _RAND_262[7:0];
  _RAND_263 = {1{`RANDOM}};
  lineBuffer_256 = _RAND_263[7:0];
  _RAND_264 = {1{`RANDOM}};
  lineBuffer_257 = _RAND_264[7:0];
  _RAND_265 = {1{`RANDOM}};
  lineBuffer_258 = _RAND_265[7:0];
  _RAND_266 = {1{`RANDOM}};
  lineBuffer_259 = _RAND_266[7:0];
  _RAND_267 = {1{`RANDOM}};
  lineBuffer_260 = _RAND_267[7:0];
  _RAND_268 = {1{`RANDOM}};
  lineBuffer_261 = _RAND_268[7:0];
  _RAND_269 = {1{`RANDOM}};
  lineBuffer_262 = _RAND_269[7:0];
  _RAND_270 = {1{`RANDOM}};
  lineBuffer_263 = _RAND_270[7:0];
  _RAND_271 = {1{`RANDOM}};
  lineBuffer_264 = _RAND_271[7:0];
  _RAND_272 = {1{`RANDOM}};
  lineBuffer_265 = _RAND_272[7:0];
  _RAND_273 = {1{`RANDOM}};
  lineBuffer_266 = _RAND_273[7:0];
  _RAND_274 = {1{`RANDOM}};
  lineBuffer_267 = _RAND_274[7:0];
  _RAND_275 = {1{`RANDOM}};
  lineBuffer_268 = _RAND_275[7:0];
  _RAND_276 = {1{`RANDOM}};
  lineBuffer_269 = _RAND_276[7:0];
  _RAND_277 = {1{`RANDOM}};
  lineBuffer_270 = _RAND_277[7:0];
  _RAND_278 = {1{`RANDOM}};
  lineBuffer_271 = _RAND_278[7:0];
  _RAND_279 = {1{`RANDOM}};
  lineBuffer_272 = _RAND_279[7:0];
  _RAND_280 = {1{`RANDOM}};
  lineBuffer_273 = _RAND_280[7:0];
  _RAND_281 = {1{`RANDOM}};
  lineBuffer_274 = _RAND_281[7:0];
  _RAND_282 = {1{`RANDOM}};
  lineBuffer_275 = _RAND_282[7:0];
  _RAND_283 = {1{`RANDOM}};
  lineBuffer_276 = _RAND_283[7:0];
  _RAND_284 = {1{`RANDOM}};
  lineBuffer_277 = _RAND_284[7:0];
  _RAND_285 = {1{`RANDOM}};
  lineBuffer_278 = _RAND_285[7:0];
  _RAND_286 = {1{`RANDOM}};
  lineBuffer_279 = _RAND_286[7:0];
  _RAND_287 = {1{`RANDOM}};
  lineBuffer_280 = _RAND_287[7:0];
  _RAND_288 = {1{`RANDOM}};
  lineBuffer_281 = _RAND_288[7:0];
  _RAND_289 = {1{`RANDOM}};
  lineBuffer_282 = _RAND_289[7:0];
  _RAND_290 = {1{`RANDOM}};
  lineBuffer_283 = _RAND_290[7:0];
  _RAND_291 = {1{`RANDOM}};
  lineBuffer_284 = _RAND_291[7:0];
  _RAND_292 = {1{`RANDOM}};
  lineBuffer_285 = _RAND_292[7:0];
  _RAND_293 = {1{`RANDOM}};
  lineBuffer_286 = _RAND_293[7:0];
  _RAND_294 = {1{`RANDOM}};
  lineBuffer_287 = _RAND_294[7:0];
  _RAND_295 = {1{`RANDOM}};
  lineBuffer_288 = _RAND_295[7:0];
  _RAND_296 = {1{`RANDOM}};
  lineBuffer_289 = _RAND_296[7:0];
  _RAND_297 = {1{`RANDOM}};
  lineBuffer_290 = _RAND_297[7:0];
  _RAND_298 = {1{`RANDOM}};
  lineBuffer_291 = _RAND_298[7:0];
  _RAND_299 = {1{`RANDOM}};
  lineBuffer_292 = _RAND_299[7:0];
  _RAND_300 = {1{`RANDOM}};
  lineBuffer_293 = _RAND_300[7:0];
  _RAND_301 = {1{`RANDOM}};
  lineBuffer_294 = _RAND_301[7:0];
  _RAND_302 = {1{`RANDOM}};
  lineBuffer_295 = _RAND_302[7:0];
  _RAND_303 = {1{`RANDOM}};
  lineBuffer_296 = _RAND_303[7:0];
  _RAND_304 = {1{`RANDOM}};
  lineBuffer_297 = _RAND_304[7:0];
  _RAND_305 = {1{`RANDOM}};
  lineBuffer_298 = _RAND_305[7:0];
  _RAND_306 = {1{`RANDOM}};
  lineBuffer_299 = _RAND_306[7:0];
  _RAND_307 = {1{`RANDOM}};
  lineBuffer_300 = _RAND_307[7:0];
  _RAND_308 = {1{`RANDOM}};
  lineBuffer_301 = _RAND_308[7:0];
  _RAND_309 = {1{`RANDOM}};
  lineBuffer_302 = _RAND_309[7:0];
  _RAND_310 = {1{`RANDOM}};
  lineBuffer_303 = _RAND_310[7:0];
  _RAND_311 = {1{`RANDOM}};
  lineBuffer_304 = _RAND_311[7:0];
  _RAND_312 = {1{`RANDOM}};
  lineBuffer_305 = _RAND_312[7:0];
  _RAND_313 = {1{`RANDOM}};
  lineBuffer_306 = _RAND_313[7:0];
  _RAND_314 = {1{`RANDOM}};
  lineBuffer_307 = _RAND_314[7:0];
  _RAND_315 = {1{`RANDOM}};
  lineBuffer_308 = _RAND_315[7:0];
  _RAND_316 = {1{`RANDOM}};
  lineBuffer_309 = _RAND_316[7:0];
  _RAND_317 = {1{`RANDOM}};
  lineBuffer_310 = _RAND_317[7:0];
  _RAND_318 = {1{`RANDOM}};
  lineBuffer_311 = _RAND_318[7:0];
  _RAND_319 = {1{`RANDOM}};
  lineBuffer_312 = _RAND_319[7:0];
  _RAND_320 = {1{`RANDOM}};
  lineBuffer_313 = _RAND_320[7:0];
  _RAND_321 = {1{`RANDOM}};
  lineBuffer_314 = _RAND_321[7:0];
  _RAND_322 = {1{`RANDOM}};
  lineBuffer_315 = _RAND_322[7:0];
  _RAND_323 = {1{`RANDOM}};
  lineBuffer_316 = _RAND_323[7:0];
  _RAND_324 = {1{`RANDOM}};
  lineBuffer_317 = _RAND_324[7:0];
  _RAND_325 = {1{`RANDOM}};
  lineBuffer_318 = _RAND_325[7:0];
  _RAND_326 = {1{`RANDOM}};
  lineBuffer_319 = _RAND_326[7:0];
  _RAND_327 = {1{`RANDOM}};
  lineBuffer_320 = _RAND_327[7:0];
  _RAND_328 = {1{`RANDOM}};
  lineBuffer_321 = _RAND_328[7:0];
  _RAND_329 = {1{`RANDOM}};
  lineBuffer_322 = _RAND_329[7:0];
  _RAND_330 = {1{`RANDOM}};
  lineBuffer_323 = _RAND_330[7:0];
  _RAND_331 = {1{`RANDOM}};
  lineBuffer_324 = _RAND_331[7:0];
  _RAND_332 = {1{`RANDOM}};
  lineBuffer_325 = _RAND_332[7:0];
  _RAND_333 = {1{`RANDOM}};
  lineBuffer_326 = _RAND_333[7:0];
  _RAND_334 = {1{`RANDOM}};
  lineBuffer_327 = _RAND_334[7:0];
  _RAND_335 = {1{`RANDOM}};
  lineBuffer_328 = _RAND_335[7:0];
  _RAND_336 = {1{`RANDOM}};
  lineBuffer_329 = _RAND_336[7:0];
  _RAND_337 = {1{`RANDOM}};
  lineBuffer_330 = _RAND_337[7:0];
  _RAND_338 = {1{`RANDOM}};
  lineBuffer_331 = _RAND_338[7:0];
  _RAND_339 = {1{`RANDOM}};
  lineBuffer_332 = _RAND_339[7:0];
  _RAND_340 = {1{`RANDOM}};
  lineBuffer_333 = _RAND_340[7:0];
  _RAND_341 = {1{`RANDOM}};
  lineBuffer_334 = _RAND_341[7:0];
  _RAND_342 = {1{`RANDOM}};
  lineBuffer_335 = _RAND_342[7:0];
  _RAND_343 = {1{`RANDOM}};
  lineBuffer_336 = _RAND_343[7:0];
  _RAND_344 = {1{`RANDOM}};
  lineBuffer_337 = _RAND_344[7:0];
  _RAND_345 = {1{`RANDOM}};
  lineBuffer_338 = _RAND_345[7:0];
  _RAND_346 = {1{`RANDOM}};
  lineBuffer_339 = _RAND_346[7:0];
  _RAND_347 = {1{`RANDOM}};
  lineBuffer_340 = _RAND_347[7:0];
  _RAND_348 = {1{`RANDOM}};
  lineBuffer_341 = _RAND_348[7:0];
  _RAND_349 = {1{`RANDOM}};
  lineBuffer_342 = _RAND_349[7:0];
  _RAND_350 = {1{`RANDOM}};
  lineBuffer_343 = _RAND_350[7:0];
  _RAND_351 = {1{`RANDOM}};
  lineBuffer_344 = _RAND_351[7:0];
  _RAND_352 = {1{`RANDOM}};
  lineBuffer_345 = _RAND_352[7:0];
  _RAND_353 = {1{`RANDOM}};
  lineBuffer_346 = _RAND_353[7:0];
  _RAND_354 = {1{`RANDOM}};
  lineBuffer_347 = _RAND_354[7:0];
  _RAND_355 = {1{`RANDOM}};
  lineBuffer_348 = _RAND_355[7:0];
  _RAND_356 = {1{`RANDOM}};
  lineBuffer_349 = _RAND_356[7:0];
  _RAND_357 = {1{`RANDOM}};
  lineBuffer_350 = _RAND_357[7:0];
  _RAND_358 = {1{`RANDOM}};
  lineBuffer_351 = _RAND_358[7:0];
  _RAND_359 = {1{`RANDOM}};
  lineBuffer_352 = _RAND_359[7:0];
  _RAND_360 = {1{`RANDOM}};
  lineBuffer_353 = _RAND_360[7:0];
  _RAND_361 = {1{`RANDOM}};
  lineBuffer_354 = _RAND_361[7:0];
  _RAND_362 = {1{`RANDOM}};
  lineBuffer_355 = _RAND_362[7:0];
  _RAND_363 = {1{`RANDOM}};
  lineBuffer_356 = _RAND_363[7:0];
  _RAND_364 = {1{`RANDOM}};
  lineBuffer_357 = _RAND_364[7:0];
  _RAND_365 = {1{`RANDOM}};
  lineBuffer_358 = _RAND_365[7:0];
  _RAND_366 = {1{`RANDOM}};
  lineBuffer_359 = _RAND_366[7:0];
  _RAND_367 = {1{`RANDOM}};
  lineBuffer_360 = _RAND_367[7:0];
  _RAND_368 = {1{`RANDOM}};
  lineBuffer_361 = _RAND_368[7:0];
  _RAND_369 = {1{`RANDOM}};
  lineBuffer_362 = _RAND_369[7:0];
  _RAND_370 = {1{`RANDOM}};
  lineBuffer_363 = _RAND_370[7:0];
  _RAND_371 = {1{`RANDOM}};
  lineBuffer_364 = _RAND_371[7:0];
  _RAND_372 = {1{`RANDOM}};
  lineBuffer_365 = _RAND_372[7:0];
  _RAND_373 = {1{`RANDOM}};
  lineBuffer_366 = _RAND_373[7:0];
  _RAND_374 = {1{`RANDOM}};
  lineBuffer_367 = _RAND_374[7:0];
  _RAND_375 = {1{`RANDOM}};
  lineBuffer_368 = _RAND_375[7:0];
  _RAND_376 = {1{`RANDOM}};
  lineBuffer_369 = _RAND_376[7:0];
  _RAND_377 = {1{`RANDOM}};
  lineBuffer_370 = _RAND_377[7:0];
  _RAND_378 = {1{`RANDOM}};
  lineBuffer_371 = _RAND_378[7:0];
  _RAND_379 = {1{`RANDOM}};
  lineBuffer_372 = _RAND_379[7:0];
  _RAND_380 = {1{`RANDOM}};
  lineBuffer_373 = _RAND_380[7:0];
  _RAND_381 = {1{`RANDOM}};
  lineBuffer_374 = _RAND_381[7:0];
  _RAND_382 = {1{`RANDOM}};
  lineBuffer_375 = _RAND_382[7:0];
  _RAND_383 = {1{`RANDOM}};
  lineBuffer_376 = _RAND_383[7:0];
  _RAND_384 = {1{`RANDOM}};
  lineBuffer_377 = _RAND_384[7:0];
  _RAND_385 = {1{`RANDOM}};
  lineBuffer_378 = _RAND_385[7:0];
  _RAND_386 = {1{`RANDOM}};
  lineBuffer_379 = _RAND_386[7:0];
  _RAND_387 = {1{`RANDOM}};
  lineBuffer_380 = _RAND_387[7:0];
  _RAND_388 = {1{`RANDOM}};
  lineBuffer_381 = _RAND_388[7:0];
  _RAND_389 = {1{`RANDOM}};
  lineBuffer_382 = _RAND_389[7:0];
  _RAND_390 = {1{`RANDOM}};
  lineBuffer_383 = _RAND_390[7:0];
  _RAND_391 = {1{`RANDOM}};
  lineBuffer_384 = _RAND_391[7:0];
  _RAND_392 = {1{`RANDOM}};
  lineBuffer_385 = _RAND_392[7:0];
  _RAND_393 = {1{`RANDOM}};
  lineBuffer_386 = _RAND_393[7:0];
  _RAND_394 = {1{`RANDOM}};
  lineBuffer_387 = _RAND_394[7:0];
  _RAND_395 = {1{`RANDOM}};
  lineBuffer_388 = _RAND_395[7:0];
  _RAND_396 = {1{`RANDOM}};
  lineBuffer_389 = _RAND_396[7:0];
  _RAND_397 = {1{`RANDOM}};
  lineBuffer_390 = _RAND_397[7:0];
  _RAND_398 = {1{`RANDOM}};
  lineBuffer_391 = _RAND_398[7:0];
  _RAND_399 = {1{`RANDOM}};
  lineBuffer_392 = _RAND_399[7:0];
  _RAND_400 = {1{`RANDOM}};
  lineBuffer_393 = _RAND_400[7:0];
  _RAND_401 = {1{`RANDOM}};
  lineBuffer_394 = _RAND_401[7:0];
  _RAND_402 = {1{`RANDOM}};
  lineBuffer_395 = _RAND_402[7:0];
  _RAND_403 = {1{`RANDOM}};
  lineBuffer_396 = _RAND_403[7:0];
  _RAND_404 = {1{`RANDOM}};
  lineBuffer_397 = _RAND_404[7:0];
  _RAND_405 = {1{`RANDOM}};
  lineBuffer_398 = _RAND_405[7:0];
  _RAND_406 = {1{`RANDOM}};
  lineBuffer_399 = _RAND_406[7:0];
  _RAND_407 = {1{`RANDOM}};
  lineBuffer_400 = _RAND_407[7:0];
  _RAND_408 = {1{`RANDOM}};
  lineBuffer_401 = _RAND_408[7:0];
  _RAND_409 = {1{`RANDOM}};
  lineBuffer_402 = _RAND_409[7:0];
  _RAND_410 = {1{`RANDOM}};
  lineBuffer_403 = _RAND_410[7:0];
  _RAND_411 = {1{`RANDOM}};
  lineBuffer_404 = _RAND_411[7:0];
  _RAND_412 = {1{`RANDOM}};
  lineBuffer_405 = _RAND_412[7:0];
  _RAND_413 = {1{`RANDOM}};
  lineBuffer_406 = _RAND_413[7:0];
  _RAND_414 = {1{`RANDOM}};
  lineBuffer_407 = _RAND_414[7:0];
  _RAND_415 = {1{`RANDOM}};
  lineBuffer_408 = _RAND_415[7:0];
  _RAND_416 = {1{`RANDOM}};
  lineBuffer_409 = _RAND_416[7:0];
  _RAND_417 = {1{`RANDOM}};
  lineBuffer_410 = _RAND_417[7:0];
  _RAND_418 = {1{`RANDOM}};
  lineBuffer_411 = _RAND_418[7:0];
  _RAND_419 = {1{`RANDOM}};
  lineBuffer_412 = _RAND_419[7:0];
  _RAND_420 = {1{`RANDOM}};
  lineBuffer_413 = _RAND_420[7:0];
  _RAND_421 = {1{`RANDOM}};
  lineBuffer_414 = _RAND_421[7:0];
  _RAND_422 = {1{`RANDOM}};
  lineBuffer_415 = _RAND_422[7:0];
  _RAND_423 = {1{`RANDOM}};
  lineBuffer_416 = _RAND_423[7:0];
  _RAND_424 = {1{`RANDOM}};
  lineBuffer_417 = _RAND_424[7:0];
  _RAND_425 = {1{`RANDOM}};
  lineBuffer_418 = _RAND_425[7:0];
  _RAND_426 = {1{`RANDOM}};
  lineBuffer_419 = _RAND_426[7:0];
  _RAND_427 = {1{`RANDOM}};
  lineBuffer_420 = _RAND_427[7:0];
  _RAND_428 = {1{`RANDOM}};
  lineBuffer_421 = _RAND_428[7:0];
  _RAND_429 = {1{`RANDOM}};
  lineBuffer_422 = _RAND_429[7:0];
  _RAND_430 = {1{`RANDOM}};
  lineBuffer_423 = _RAND_430[7:0];
  _RAND_431 = {1{`RANDOM}};
  lineBuffer_424 = _RAND_431[7:0];
  _RAND_432 = {1{`RANDOM}};
  lineBuffer_425 = _RAND_432[7:0];
  _RAND_433 = {1{`RANDOM}};
  lineBuffer_426 = _RAND_433[7:0];
  _RAND_434 = {1{`RANDOM}};
  lineBuffer_427 = _RAND_434[7:0];
  _RAND_435 = {1{`RANDOM}};
  lineBuffer_428 = _RAND_435[7:0];
  _RAND_436 = {1{`RANDOM}};
  lineBuffer_429 = _RAND_436[7:0];
  _RAND_437 = {1{`RANDOM}};
  lineBuffer_430 = _RAND_437[7:0];
  _RAND_438 = {1{`RANDOM}};
  lineBuffer_431 = _RAND_438[7:0];
  _RAND_439 = {1{`RANDOM}};
  lineBuffer_432 = _RAND_439[7:0];
  _RAND_440 = {1{`RANDOM}};
  lineBuffer_433 = _RAND_440[7:0];
  _RAND_441 = {1{`RANDOM}};
  lineBuffer_434 = _RAND_441[7:0];
  _RAND_442 = {1{`RANDOM}};
  lineBuffer_435 = _RAND_442[7:0];
  _RAND_443 = {1{`RANDOM}};
  lineBuffer_436 = _RAND_443[7:0];
  _RAND_444 = {1{`RANDOM}};
  lineBuffer_437 = _RAND_444[7:0];
  _RAND_445 = {1{`RANDOM}};
  lineBuffer_438 = _RAND_445[7:0];
  _RAND_446 = {1{`RANDOM}};
  lineBuffer_439 = _RAND_446[7:0];
  _RAND_447 = {1{`RANDOM}};
  lineBuffer_440 = _RAND_447[7:0];
  _RAND_448 = {1{`RANDOM}};
  lineBuffer_441 = _RAND_448[7:0];
  _RAND_449 = {1{`RANDOM}};
  lineBuffer_442 = _RAND_449[7:0];
  _RAND_450 = {1{`RANDOM}};
  lineBuffer_443 = _RAND_450[7:0];
  _RAND_451 = {1{`RANDOM}};
  lineBuffer_444 = _RAND_451[7:0];
  _RAND_452 = {1{`RANDOM}};
  lineBuffer_445 = _RAND_452[7:0];
  _RAND_453 = {1{`RANDOM}};
  lineBuffer_446 = _RAND_453[7:0];
  _RAND_454 = {1{`RANDOM}};
  lineBuffer_447 = _RAND_454[7:0];
  _RAND_455 = {1{`RANDOM}};
  lineBuffer_448 = _RAND_455[7:0];
  _RAND_456 = {1{`RANDOM}};
  lineBuffer_449 = _RAND_456[7:0];
  _RAND_457 = {1{`RANDOM}};
  lineBuffer_450 = _RAND_457[7:0];
  _RAND_458 = {1{`RANDOM}};
  lineBuffer_451 = _RAND_458[7:0];
  _RAND_459 = {1{`RANDOM}};
  lineBuffer_452 = _RAND_459[7:0];
  _RAND_460 = {1{`RANDOM}};
  lineBuffer_453 = _RAND_460[7:0];
  _RAND_461 = {1{`RANDOM}};
  lineBuffer_454 = _RAND_461[7:0];
  _RAND_462 = {1{`RANDOM}};
  lineBuffer_455 = _RAND_462[7:0];
  _RAND_463 = {1{`RANDOM}};
  lineBuffer_456 = _RAND_463[7:0];
  _RAND_464 = {1{`RANDOM}};
  lineBuffer_457 = _RAND_464[7:0];
  _RAND_465 = {1{`RANDOM}};
  lineBuffer_458 = _RAND_465[7:0];
  _RAND_466 = {1{`RANDOM}};
  lineBuffer_459 = _RAND_466[7:0];
  _RAND_467 = {1{`RANDOM}};
  lineBuffer_460 = _RAND_467[7:0];
  _RAND_468 = {1{`RANDOM}};
  lineBuffer_461 = _RAND_468[7:0];
  _RAND_469 = {1{`RANDOM}};
  lineBuffer_462 = _RAND_469[7:0];
  _RAND_470 = {1{`RANDOM}};
  lineBuffer_463 = _RAND_470[7:0];
  _RAND_471 = {1{`RANDOM}};
  lineBuffer_464 = _RAND_471[7:0];
  _RAND_472 = {1{`RANDOM}};
  lineBuffer_465 = _RAND_472[7:0];
  _RAND_473 = {1{`RANDOM}};
  lineBuffer_466 = _RAND_473[7:0];
  _RAND_474 = {1{`RANDOM}};
  lineBuffer_467 = _RAND_474[7:0];
  _RAND_475 = {1{`RANDOM}};
  lineBuffer_468 = _RAND_475[7:0];
  _RAND_476 = {1{`RANDOM}};
  lineBuffer_469 = _RAND_476[7:0];
  _RAND_477 = {1{`RANDOM}};
  lineBuffer_470 = _RAND_477[7:0];
  _RAND_478 = {1{`RANDOM}};
  lineBuffer_471 = _RAND_478[7:0];
  _RAND_479 = {1{`RANDOM}};
  lineBuffer_472 = _RAND_479[7:0];
  _RAND_480 = {1{`RANDOM}};
  lineBuffer_473 = _RAND_480[7:0];
  _RAND_481 = {1{`RANDOM}};
  lineBuffer_474 = _RAND_481[7:0];
  _RAND_482 = {1{`RANDOM}};
  lineBuffer_475 = _RAND_482[7:0];
  _RAND_483 = {1{`RANDOM}};
  lineBuffer_476 = _RAND_483[7:0];
  _RAND_484 = {1{`RANDOM}};
  lineBuffer_477 = _RAND_484[7:0];
  _RAND_485 = {1{`RANDOM}};
  lineBuffer_478 = _RAND_485[7:0];
  _RAND_486 = {1{`RANDOM}};
  lineBuffer_479 = _RAND_486[7:0];
  _RAND_487 = {1{`RANDOM}};
  lineBuffer_480 = _RAND_487[7:0];
  _RAND_488 = {1{`RANDOM}};
  lineBuffer_481 = _RAND_488[7:0];
  _RAND_489 = {1{`RANDOM}};
  lineBuffer_482 = _RAND_489[7:0];
  _RAND_490 = {1{`RANDOM}};
  lineBuffer_483 = _RAND_490[7:0];
  _RAND_491 = {1{`RANDOM}};
  lineBuffer_484 = _RAND_491[7:0];
  _RAND_492 = {1{`RANDOM}};
  lineBuffer_485 = _RAND_492[7:0];
  _RAND_493 = {1{`RANDOM}};
  lineBuffer_486 = _RAND_493[7:0];
  _RAND_494 = {1{`RANDOM}};
  lineBuffer_487 = _RAND_494[7:0];
  _RAND_495 = {1{`RANDOM}};
  lineBuffer_488 = _RAND_495[7:0];
  _RAND_496 = {1{`RANDOM}};
  lineBuffer_489 = _RAND_496[7:0];
  _RAND_497 = {1{`RANDOM}};
  lineBuffer_490 = _RAND_497[7:0];
  _RAND_498 = {1{`RANDOM}};
  lineBuffer_491 = _RAND_498[7:0];
  _RAND_499 = {1{`RANDOM}};
  lineBuffer_492 = _RAND_499[7:0];
  _RAND_500 = {1{`RANDOM}};
  lineBuffer_493 = _RAND_500[7:0];
  _RAND_501 = {1{`RANDOM}};
  lineBuffer_494 = _RAND_501[7:0];
  _RAND_502 = {1{`RANDOM}};
  lineBuffer_495 = _RAND_502[7:0];
  _RAND_503 = {1{`RANDOM}};
  lineBuffer_496 = _RAND_503[7:0];
  _RAND_504 = {1{`RANDOM}};
  lineBuffer_497 = _RAND_504[7:0];
  _RAND_505 = {1{`RANDOM}};
  lineBuffer_498 = _RAND_505[7:0];
  _RAND_506 = {1{`RANDOM}};
  lineBuffer_499 = _RAND_506[7:0];
  _RAND_507 = {1{`RANDOM}};
  lineBuffer_500 = _RAND_507[7:0];
  _RAND_508 = {1{`RANDOM}};
  lineBuffer_501 = _RAND_508[7:0];
  _RAND_509 = {1{`RANDOM}};
  lineBuffer_502 = _RAND_509[7:0];
  _RAND_510 = {1{`RANDOM}};
  lineBuffer_503 = _RAND_510[7:0];
  _RAND_511 = {1{`RANDOM}};
  lineBuffer_504 = _RAND_511[7:0];
  _RAND_512 = {1{`RANDOM}};
  lineBuffer_505 = _RAND_512[7:0];
  _RAND_513 = {1{`RANDOM}};
  lineBuffer_506 = _RAND_513[7:0];
  _RAND_514 = {1{`RANDOM}};
  lineBuffer_507 = _RAND_514[7:0];
  _RAND_515 = {1{`RANDOM}};
  lineBuffer_508 = _RAND_515[7:0];
  _RAND_516 = {1{`RANDOM}};
  lineBuffer_509 = _RAND_516[7:0];
  _RAND_517 = {1{`RANDOM}};
  lineBuffer_510 = _RAND_517[7:0];
  _RAND_518 = {1{`RANDOM}};
  lineBuffer_511 = _RAND_518[7:0];
  _RAND_519 = {1{`RANDOM}};
  lineBuffer_512 = _RAND_519[7:0];
  _RAND_520 = {1{`RANDOM}};
  lineBuffer_513 = _RAND_520[7:0];
  _RAND_521 = {1{`RANDOM}};
  lineBuffer_514 = _RAND_521[7:0];
  _RAND_522 = {1{`RANDOM}};
  lineBuffer_515 = _RAND_522[7:0];
  _RAND_523 = {1{`RANDOM}};
  lineBuffer_516 = _RAND_523[7:0];
  _RAND_524 = {1{`RANDOM}};
  lineBuffer_517 = _RAND_524[7:0];
  _RAND_525 = {1{`RANDOM}};
  lineBuffer_518 = _RAND_525[7:0];
  _RAND_526 = {1{`RANDOM}};
  lineBuffer_519 = _RAND_526[7:0];
  _RAND_527 = {1{`RANDOM}};
  lineBuffer_520 = _RAND_527[7:0];
  _RAND_528 = {1{`RANDOM}};
  lineBuffer_521 = _RAND_528[7:0];
  _RAND_529 = {1{`RANDOM}};
  lineBuffer_522 = _RAND_529[7:0];
  _RAND_530 = {1{`RANDOM}};
  lineBuffer_523 = _RAND_530[7:0];
  _RAND_531 = {1{`RANDOM}};
  lineBuffer_524 = _RAND_531[7:0];
  _RAND_532 = {1{`RANDOM}};
  lineBuffer_525 = _RAND_532[7:0];
  _RAND_533 = {1{`RANDOM}};
  lineBuffer_526 = _RAND_533[7:0];
  _RAND_534 = {1{`RANDOM}};
  lineBuffer_527 = _RAND_534[7:0];
  _RAND_535 = {1{`RANDOM}};
  lineBuffer_528 = _RAND_535[7:0];
  _RAND_536 = {1{`RANDOM}};
  lineBuffer_529 = _RAND_536[7:0];
  _RAND_537 = {1{`RANDOM}};
  lineBuffer_530 = _RAND_537[7:0];
  _RAND_538 = {1{`RANDOM}};
  lineBuffer_531 = _RAND_538[7:0];
  _RAND_539 = {1{`RANDOM}};
  lineBuffer_532 = _RAND_539[7:0];
  _RAND_540 = {1{`RANDOM}};
  lineBuffer_533 = _RAND_540[7:0];
  _RAND_541 = {1{`RANDOM}};
  lineBuffer_534 = _RAND_541[7:0];
  _RAND_542 = {1{`RANDOM}};
  lineBuffer_535 = _RAND_542[7:0];
  _RAND_543 = {1{`RANDOM}};
  lineBuffer_536 = _RAND_543[7:0];
  _RAND_544 = {1{`RANDOM}};
  lineBuffer_537 = _RAND_544[7:0];
  _RAND_545 = {1{`RANDOM}};
  lineBuffer_538 = _RAND_545[7:0];
  _RAND_546 = {1{`RANDOM}};
  lineBuffer_539 = _RAND_546[7:0];
  _RAND_547 = {1{`RANDOM}};
  lineBuffer_540 = _RAND_547[7:0];
  _RAND_548 = {1{`RANDOM}};
  lineBuffer_541 = _RAND_548[7:0];
  _RAND_549 = {1{`RANDOM}};
  lineBuffer_542 = _RAND_549[7:0];
  _RAND_550 = {1{`RANDOM}};
  lineBuffer_543 = _RAND_550[7:0];
  _RAND_551 = {1{`RANDOM}};
  lineBuffer_544 = _RAND_551[7:0];
  _RAND_552 = {1{`RANDOM}};
  lineBuffer_545 = _RAND_552[7:0];
  _RAND_553 = {1{`RANDOM}};
  lineBuffer_546 = _RAND_553[7:0];
  _RAND_554 = {1{`RANDOM}};
  lineBuffer_547 = _RAND_554[7:0];
  _RAND_555 = {1{`RANDOM}};
  lineBuffer_548 = _RAND_555[7:0];
  _RAND_556 = {1{`RANDOM}};
  lineBuffer_549 = _RAND_556[7:0];
  _RAND_557 = {1{`RANDOM}};
  lineBuffer_550 = _RAND_557[7:0];
  _RAND_558 = {1{`RANDOM}};
  lineBuffer_551 = _RAND_558[7:0];
  _RAND_559 = {1{`RANDOM}};
  lineBuffer_552 = _RAND_559[7:0];
  _RAND_560 = {1{`RANDOM}};
  lineBuffer_553 = _RAND_560[7:0];
  _RAND_561 = {1{`RANDOM}};
  lineBuffer_554 = _RAND_561[7:0];
  _RAND_562 = {1{`RANDOM}};
  lineBuffer_555 = _RAND_562[7:0];
  _RAND_563 = {1{`RANDOM}};
  lineBuffer_556 = _RAND_563[7:0];
  _RAND_564 = {1{`RANDOM}};
  lineBuffer_557 = _RAND_564[7:0];
  _RAND_565 = {1{`RANDOM}};
  lineBuffer_558 = _RAND_565[7:0];
  _RAND_566 = {1{`RANDOM}};
  lineBuffer_559 = _RAND_566[7:0];
  _RAND_567 = {1{`RANDOM}};
  lineBuffer_560 = _RAND_567[7:0];
  _RAND_568 = {1{`RANDOM}};
  lineBuffer_561 = _RAND_568[7:0];
  _RAND_569 = {1{`RANDOM}};
  lineBuffer_562 = _RAND_569[7:0];
  _RAND_570 = {1{`RANDOM}};
  lineBuffer_563 = _RAND_570[7:0];
  _RAND_571 = {1{`RANDOM}};
  lineBuffer_564 = _RAND_571[7:0];
  _RAND_572 = {1{`RANDOM}};
  lineBuffer_565 = _RAND_572[7:0];
  _RAND_573 = {1{`RANDOM}};
  lineBuffer_566 = _RAND_573[7:0];
  _RAND_574 = {1{`RANDOM}};
  lineBuffer_567 = _RAND_574[7:0];
  _RAND_575 = {1{`RANDOM}};
  lineBuffer_568 = _RAND_575[7:0];
  _RAND_576 = {1{`RANDOM}};
  lineBuffer_569 = _RAND_576[7:0];
  _RAND_577 = {1{`RANDOM}};
  lineBuffer_570 = _RAND_577[7:0];
  _RAND_578 = {1{`RANDOM}};
  lineBuffer_571 = _RAND_578[7:0];
  _RAND_579 = {1{`RANDOM}};
  lineBuffer_572 = _RAND_579[7:0];
  _RAND_580 = {1{`RANDOM}};
  lineBuffer_573 = _RAND_580[7:0];
  _RAND_581 = {1{`RANDOM}};
  lineBuffer_574 = _RAND_581[7:0];
  _RAND_582 = {1{`RANDOM}};
  lineBuffer_575 = _RAND_582[7:0];
  _RAND_583 = {1{`RANDOM}};
  lineBuffer_576 = _RAND_583[7:0];
  _RAND_584 = {1{`RANDOM}};
  lineBuffer_577 = _RAND_584[7:0];
  _RAND_585 = {1{`RANDOM}};
  lineBuffer_578 = _RAND_585[7:0];
  _RAND_586 = {1{`RANDOM}};
  lineBuffer_579 = _RAND_586[7:0];
  _RAND_587 = {1{`RANDOM}};
  lineBuffer_580 = _RAND_587[7:0];
  _RAND_588 = {1{`RANDOM}};
  lineBuffer_581 = _RAND_588[7:0];
  _RAND_589 = {1{`RANDOM}};
  lineBuffer_582 = _RAND_589[7:0];
  _RAND_590 = {1{`RANDOM}};
  lineBuffer_583 = _RAND_590[7:0];
  _RAND_591 = {1{`RANDOM}};
  lineBuffer_584 = _RAND_591[7:0];
  _RAND_592 = {1{`RANDOM}};
  lineBuffer_585 = _RAND_592[7:0];
  _RAND_593 = {1{`RANDOM}};
  lineBuffer_586 = _RAND_593[7:0];
  _RAND_594 = {1{`RANDOM}};
  lineBuffer_587 = _RAND_594[7:0];
  _RAND_595 = {1{`RANDOM}};
  lineBuffer_588 = _RAND_595[7:0];
  _RAND_596 = {1{`RANDOM}};
  lineBuffer_589 = _RAND_596[7:0];
  _RAND_597 = {1{`RANDOM}};
  lineBuffer_590 = _RAND_597[7:0];
  _RAND_598 = {1{`RANDOM}};
  lineBuffer_591 = _RAND_598[7:0];
  _RAND_599 = {1{`RANDOM}};
  lineBuffer_592 = _RAND_599[7:0];
  _RAND_600 = {1{`RANDOM}};
  lineBuffer_593 = _RAND_600[7:0];
  _RAND_601 = {1{`RANDOM}};
  lineBuffer_594 = _RAND_601[7:0];
  _RAND_602 = {1{`RANDOM}};
  lineBuffer_595 = _RAND_602[7:0];
  _RAND_603 = {1{`RANDOM}};
  lineBuffer_596 = _RAND_603[7:0];
  _RAND_604 = {1{`RANDOM}};
  lineBuffer_597 = _RAND_604[7:0];
  _RAND_605 = {1{`RANDOM}};
  lineBuffer_598 = _RAND_605[7:0];
  _RAND_606 = {1{`RANDOM}};
  lineBuffer_599 = _RAND_606[7:0];
  _RAND_607 = {1{`RANDOM}};
  lineBuffer_600 = _RAND_607[7:0];
  _RAND_608 = {1{`RANDOM}};
  lineBuffer_601 = _RAND_608[7:0];
  _RAND_609 = {1{`RANDOM}};
  lineBuffer_602 = _RAND_609[7:0];
  _RAND_610 = {1{`RANDOM}};
  lineBuffer_603 = _RAND_610[7:0];
  _RAND_611 = {1{`RANDOM}};
  lineBuffer_604 = _RAND_611[7:0];
  _RAND_612 = {1{`RANDOM}};
  lineBuffer_605 = _RAND_612[7:0];
  _RAND_613 = {1{`RANDOM}};
  lineBuffer_606 = _RAND_613[7:0];
  _RAND_614 = {1{`RANDOM}};
  lineBuffer_607 = _RAND_614[7:0];
  _RAND_615 = {1{`RANDOM}};
  lineBuffer_608 = _RAND_615[7:0];
  _RAND_616 = {1{`RANDOM}};
  lineBuffer_609 = _RAND_616[7:0];
  _RAND_617 = {1{`RANDOM}};
  lineBuffer_610 = _RAND_617[7:0];
  _RAND_618 = {1{`RANDOM}};
  lineBuffer_611 = _RAND_618[7:0];
  _RAND_619 = {1{`RANDOM}};
  lineBuffer_612 = _RAND_619[7:0];
  _RAND_620 = {1{`RANDOM}};
  lineBuffer_613 = _RAND_620[7:0];
  _RAND_621 = {1{`RANDOM}};
  lineBuffer_614 = _RAND_621[7:0];
  _RAND_622 = {1{`RANDOM}};
  lineBuffer_615 = _RAND_622[7:0];
  _RAND_623 = {1{`RANDOM}};
  lineBuffer_616 = _RAND_623[7:0];
  _RAND_624 = {1{`RANDOM}};
  lineBuffer_617 = _RAND_624[7:0];
  _RAND_625 = {1{`RANDOM}};
  lineBuffer_618 = _RAND_625[7:0];
  _RAND_626 = {1{`RANDOM}};
  lineBuffer_619 = _RAND_626[7:0];
  _RAND_627 = {1{`RANDOM}};
  lineBuffer_620 = _RAND_627[7:0];
  _RAND_628 = {1{`RANDOM}};
  lineBuffer_621 = _RAND_628[7:0];
  _RAND_629 = {1{`RANDOM}};
  lineBuffer_622 = _RAND_629[7:0];
  _RAND_630 = {1{`RANDOM}};
  lineBuffer_623 = _RAND_630[7:0];
  _RAND_631 = {1{`RANDOM}};
  lineBuffer_624 = _RAND_631[7:0];
  _RAND_632 = {1{`RANDOM}};
  lineBuffer_625 = _RAND_632[7:0];
  _RAND_633 = {1{`RANDOM}};
  lineBuffer_626 = _RAND_633[7:0];
  _RAND_634 = {1{`RANDOM}};
  lineBuffer_627 = _RAND_634[7:0];
  _RAND_635 = {1{`RANDOM}};
  lineBuffer_628 = _RAND_635[7:0];
  _RAND_636 = {1{`RANDOM}};
  lineBuffer_629 = _RAND_636[7:0];
  _RAND_637 = {1{`RANDOM}};
  lineBuffer_630 = _RAND_637[7:0];
  _RAND_638 = {1{`RANDOM}};
  lineBuffer_631 = _RAND_638[7:0];
  _RAND_639 = {1{`RANDOM}};
  lineBuffer_632 = _RAND_639[7:0];
  _RAND_640 = {1{`RANDOM}};
  lineBuffer_633 = _RAND_640[7:0];
  _RAND_641 = {1{`RANDOM}};
  lineBuffer_634 = _RAND_641[7:0];
  _RAND_642 = {1{`RANDOM}};
  lineBuffer_635 = _RAND_642[7:0];
  _RAND_643 = {1{`RANDOM}};
  lineBuffer_636 = _RAND_643[7:0];
  _RAND_644 = {1{`RANDOM}};
  lineBuffer_637 = _RAND_644[7:0];
  _RAND_645 = {1{`RANDOM}};
  lineBuffer_638 = _RAND_645[7:0];
  _RAND_646 = {1{`RANDOM}};
  lineBuffer_639 = _RAND_646[7:0];
  _RAND_647 = {1{`RANDOM}};
  lineBuffer_640 = _RAND_647[7:0];
  _RAND_648 = {1{`RANDOM}};
  lineBuffer_641 = _RAND_648[7:0];
  _RAND_649 = {1{`RANDOM}};
  lineBuffer_642 = _RAND_649[7:0];
  _RAND_650 = {1{`RANDOM}};
  lineBuffer_643 = _RAND_650[7:0];
  _RAND_651 = {1{`RANDOM}};
  lineBuffer_644 = _RAND_651[7:0];
  _RAND_652 = {1{`RANDOM}};
  lineBuffer_645 = _RAND_652[7:0];
  _RAND_653 = {1{`RANDOM}};
  lineBuffer_646 = _RAND_653[7:0];
  _RAND_654 = {1{`RANDOM}};
  lineBuffer_647 = _RAND_654[7:0];
  _RAND_655 = {1{`RANDOM}};
  lineBuffer_648 = _RAND_655[7:0];
  _RAND_656 = {1{`RANDOM}};
  lineBuffer_649 = _RAND_656[7:0];
  _RAND_657 = {1{`RANDOM}};
  lineBuffer_650 = _RAND_657[7:0];
  _RAND_658 = {1{`RANDOM}};
  lineBuffer_651 = _RAND_658[7:0];
  _RAND_659 = {1{`RANDOM}};
  lineBuffer_652 = _RAND_659[7:0];
  _RAND_660 = {1{`RANDOM}};
  lineBuffer_653 = _RAND_660[7:0];
  _RAND_661 = {1{`RANDOM}};
  lineBuffer_654 = _RAND_661[7:0];
  _RAND_662 = {1{`RANDOM}};
  lineBuffer_655 = _RAND_662[7:0];
  _RAND_663 = {1{`RANDOM}};
  lineBuffer_656 = _RAND_663[7:0];
  _RAND_664 = {1{`RANDOM}};
  lineBuffer_657 = _RAND_664[7:0];
  _RAND_665 = {1{`RANDOM}};
  lineBuffer_658 = _RAND_665[7:0];
  _RAND_666 = {1{`RANDOM}};
  lineBuffer_659 = _RAND_666[7:0];
  _RAND_667 = {1{`RANDOM}};
  lineBuffer_660 = _RAND_667[7:0];
  _RAND_668 = {1{`RANDOM}};
  lineBuffer_661 = _RAND_668[7:0];
  _RAND_669 = {1{`RANDOM}};
  lineBuffer_662 = _RAND_669[7:0];
  _RAND_670 = {1{`RANDOM}};
  lineBuffer_663 = _RAND_670[7:0];
  _RAND_671 = {1{`RANDOM}};
  lineBuffer_664 = _RAND_671[7:0];
  _RAND_672 = {1{`RANDOM}};
  lineBuffer_665 = _RAND_672[7:0];
  _RAND_673 = {1{`RANDOM}};
  lineBuffer_666 = _RAND_673[7:0];
  _RAND_674 = {1{`RANDOM}};
  lineBuffer_667 = _RAND_674[7:0];
  _RAND_675 = {1{`RANDOM}};
  lineBuffer_668 = _RAND_675[7:0];
  _RAND_676 = {1{`RANDOM}};
  lineBuffer_669 = _RAND_676[7:0];
  _RAND_677 = {1{`RANDOM}};
  lineBuffer_670 = _RAND_677[7:0];
  _RAND_678 = {1{`RANDOM}};
  lineBuffer_671 = _RAND_678[7:0];
  _RAND_679 = {1{`RANDOM}};
  lineBuffer_672 = _RAND_679[7:0];
  _RAND_680 = {1{`RANDOM}};
  lineBuffer_673 = _RAND_680[7:0];
  _RAND_681 = {1{`RANDOM}};
  lineBuffer_674 = _RAND_681[7:0];
  _RAND_682 = {1{`RANDOM}};
  lineBuffer_675 = _RAND_682[7:0];
  _RAND_683 = {1{`RANDOM}};
  lineBuffer_676 = _RAND_683[7:0];
  _RAND_684 = {1{`RANDOM}};
  lineBuffer_677 = _RAND_684[7:0];
  _RAND_685 = {1{`RANDOM}};
  lineBuffer_678 = _RAND_685[7:0];
  _RAND_686 = {1{`RANDOM}};
  lineBuffer_679 = _RAND_686[7:0];
  _RAND_687 = {1{`RANDOM}};
  lineBuffer_680 = _RAND_687[7:0];
  _RAND_688 = {1{`RANDOM}};
  lineBuffer_681 = _RAND_688[7:0];
  _RAND_689 = {1{`RANDOM}};
  lineBuffer_682 = _RAND_689[7:0];
  _RAND_690 = {1{`RANDOM}};
  lineBuffer_683 = _RAND_690[7:0];
  _RAND_691 = {1{`RANDOM}};
  lineBuffer_684 = _RAND_691[7:0];
  _RAND_692 = {1{`RANDOM}};
  lineBuffer_685 = _RAND_692[7:0];
  _RAND_693 = {1{`RANDOM}};
  lineBuffer_686 = _RAND_693[7:0];
  _RAND_694 = {1{`RANDOM}};
  lineBuffer_687 = _RAND_694[7:0];
  _RAND_695 = {1{`RANDOM}};
  lineBuffer_688 = _RAND_695[7:0];
  _RAND_696 = {1{`RANDOM}};
  lineBuffer_689 = _RAND_696[7:0];
  _RAND_697 = {1{`RANDOM}};
  lineBuffer_690 = _RAND_697[7:0];
  _RAND_698 = {1{`RANDOM}};
  lineBuffer_691 = _RAND_698[7:0];
  _RAND_699 = {1{`RANDOM}};
  lineBuffer_692 = _RAND_699[7:0];
  _RAND_700 = {1{`RANDOM}};
  lineBuffer_693 = _RAND_700[7:0];
  _RAND_701 = {1{`RANDOM}};
  lineBuffer_694 = _RAND_701[7:0];
  _RAND_702 = {1{`RANDOM}};
  lineBuffer_695 = _RAND_702[7:0];
  _RAND_703 = {1{`RANDOM}};
  lineBuffer_696 = _RAND_703[7:0];
  _RAND_704 = {1{`RANDOM}};
  lineBuffer_697 = _RAND_704[7:0];
  _RAND_705 = {1{`RANDOM}};
  lineBuffer_698 = _RAND_705[7:0];
  _RAND_706 = {1{`RANDOM}};
  lineBuffer_699 = _RAND_706[7:0];
  _RAND_707 = {1{`RANDOM}};
  lineBuffer_700 = _RAND_707[7:0];
  _RAND_708 = {1{`RANDOM}};
  lineBuffer_701 = _RAND_708[7:0];
  _RAND_709 = {1{`RANDOM}};
  lineBuffer_702 = _RAND_709[7:0];
  _RAND_710 = {1{`RANDOM}};
  lineBuffer_703 = _RAND_710[7:0];
  _RAND_711 = {1{`RANDOM}};
  lineBuffer_704 = _RAND_711[7:0];
  _RAND_712 = {1{`RANDOM}};
  lineBuffer_705 = _RAND_712[7:0];
  _RAND_713 = {1{`RANDOM}};
  lineBuffer_706 = _RAND_713[7:0];
  _RAND_714 = {1{`RANDOM}};
  lineBuffer_707 = _RAND_714[7:0];
  _RAND_715 = {1{`RANDOM}};
  lineBuffer_708 = _RAND_715[7:0];
  _RAND_716 = {1{`RANDOM}};
  lineBuffer_709 = _RAND_716[7:0];
  _RAND_717 = {1{`RANDOM}};
  lineBuffer_710 = _RAND_717[7:0];
  _RAND_718 = {1{`RANDOM}};
  lineBuffer_711 = _RAND_718[7:0];
  _RAND_719 = {1{`RANDOM}};
  lineBuffer_712 = _RAND_719[7:0];
  _RAND_720 = {1{`RANDOM}};
  lineBuffer_713 = _RAND_720[7:0];
  _RAND_721 = {1{`RANDOM}};
  lineBuffer_714 = _RAND_721[7:0];
  _RAND_722 = {1{`RANDOM}};
  lineBuffer_715 = _RAND_722[7:0];
  _RAND_723 = {1{`RANDOM}};
  lineBuffer_716 = _RAND_723[7:0];
  _RAND_724 = {1{`RANDOM}};
  lineBuffer_717 = _RAND_724[7:0];
  _RAND_725 = {1{`RANDOM}};
  lineBuffer_718 = _RAND_725[7:0];
  _RAND_726 = {1{`RANDOM}};
  lineBuffer_719 = _RAND_726[7:0];
  _RAND_727 = {1{`RANDOM}};
  lineBuffer_720 = _RAND_727[7:0];
  _RAND_728 = {1{`RANDOM}};
  lineBuffer_721 = _RAND_728[7:0];
  _RAND_729 = {1{`RANDOM}};
  lineBuffer_722 = _RAND_729[7:0];
  _RAND_730 = {1{`RANDOM}};
  lineBuffer_723 = _RAND_730[7:0];
  _RAND_731 = {1{`RANDOM}};
  lineBuffer_724 = _RAND_731[7:0];
  _RAND_732 = {1{`RANDOM}};
  lineBuffer_725 = _RAND_732[7:0];
  _RAND_733 = {1{`RANDOM}};
  lineBuffer_726 = _RAND_733[7:0];
  _RAND_734 = {1{`RANDOM}};
  lineBuffer_727 = _RAND_734[7:0];
  _RAND_735 = {1{`RANDOM}};
  lineBuffer_728 = _RAND_735[7:0];
  _RAND_736 = {1{`RANDOM}};
  lineBuffer_729 = _RAND_736[7:0];
  _RAND_737 = {1{`RANDOM}};
  lineBuffer_730 = _RAND_737[7:0];
  _RAND_738 = {1{`RANDOM}};
  lineBuffer_731 = _RAND_738[7:0];
  _RAND_739 = {1{`RANDOM}};
  lineBuffer_732 = _RAND_739[7:0];
  _RAND_740 = {1{`RANDOM}};
  lineBuffer_733 = _RAND_740[7:0];
  _RAND_741 = {1{`RANDOM}};
  lineBuffer_734 = _RAND_741[7:0];
  _RAND_742 = {1{`RANDOM}};
  lineBuffer_735 = _RAND_742[7:0];
  _RAND_743 = {1{`RANDOM}};
  lineBuffer_736 = _RAND_743[7:0];
  _RAND_744 = {1{`RANDOM}};
  lineBuffer_737 = _RAND_744[7:0];
  _RAND_745 = {1{`RANDOM}};
  lineBuffer_738 = _RAND_745[7:0];
  _RAND_746 = {1{`RANDOM}};
  lineBuffer_739 = _RAND_746[7:0];
  _RAND_747 = {1{`RANDOM}};
  lineBuffer_740 = _RAND_747[7:0];
  _RAND_748 = {1{`RANDOM}};
  lineBuffer_741 = _RAND_748[7:0];
  _RAND_749 = {1{`RANDOM}};
  lineBuffer_742 = _RAND_749[7:0];
  _RAND_750 = {1{`RANDOM}};
  lineBuffer_743 = _RAND_750[7:0];
  _RAND_751 = {1{`RANDOM}};
  lineBuffer_744 = _RAND_751[7:0];
  _RAND_752 = {1{`RANDOM}};
  lineBuffer_745 = _RAND_752[7:0];
  _RAND_753 = {1{`RANDOM}};
  lineBuffer_746 = _RAND_753[7:0];
  _RAND_754 = {1{`RANDOM}};
  lineBuffer_747 = _RAND_754[7:0];
  _RAND_755 = {1{`RANDOM}};
  lineBuffer_748 = _RAND_755[7:0];
  _RAND_756 = {1{`RANDOM}};
  lineBuffer_749 = _RAND_756[7:0];
  _RAND_757 = {1{`RANDOM}};
  lineBuffer_750 = _RAND_757[7:0];
  _RAND_758 = {1{`RANDOM}};
  lineBuffer_751 = _RAND_758[7:0];
  _RAND_759 = {1{`RANDOM}};
  lineBuffer_752 = _RAND_759[7:0];
  _RAND_760 = {1{`RANDOM}};
  lineBuffer_753 = _RAND_760[7:0];
  _RAND_761 = {1{`RANDOM}};
  lineBuffer_754 = _RAND_761[7:0];
  _RAND_762 = {1{`RANDOM}};
  lineBuffer_755 = _RAND_762[7:0];
  _RAND_763 = {1{`RANDOM}};
  lineBuffer_756 = _RAND_763[7:0];
  _RAND_764 = {1{`RANDOM}};
  lineBuffer_757 = _RAND_764[7:0];
  _RAND_765 = {1{`RANDOM}};
  lineBuffer_758 = _RAND_765[7:0];
  _RAND_766 = {1{`RANDOM}};
  lineBuffer_759 = _RAND_766[7:0];
  _RAND_767 = {1{`RANDOM}};
  lineBuffer_760 = _RAND_767[7:0];
  _RAND_768 = {1{`RANDOM}};
  lineBuffer_761 = _RAND_768[7:0];
  _RAND_769 = {1{`RANDOM}};
  lineBuffer_762 = _RAND_769[7:0];
  _RAND_770 = {1{`RANDOM}};
  lineBuffer_763 = _RAND_770[7:0];
  _RAND_771 = {1{`RANDOM}};
  lineBuffer_764 = _RAND_771[7:0];
  _RAND_772 = {1{`RANDOM}};
  lineBuffer_765 = _RAND_772[7:0];
  _RAND_773 = {1{`RANDOM}};
  lineBuffer_766 = _RAND_773[7:0];
  _RAND_774 = {1{`RANDOM}};
  lineBuffer_767 = _RAND_774[7:0];
  _RAND_775 = {1{`RANDOM}};
  windowBuffer_0 = _RAND_775[15:0];
  _RAND_776 = {1{`RANDOM}};
  windowBuffer_1 = _RAND_776[15:0];
  _RAND_777 = {1{`RANDOM}};
  windowBuffer_2 = _RAND_777[15:0];
  _RAND_778 = {1{`RANDOM}};
  windowBuffer_3 = _RAND_778[15:0];
  _RAND_779 = {1{`RANDOM}};
  windowBuffer_4 = _RAND_779[15:0];
  _RAND_780 = {1{`RANDOM}};
  windowBuffer_5 = _RAND_780[15:0];
  _RAND_781 = {1{`RANDOM}};
  windowBuffer_6 = _RAND_781[15:0];
  _RAND_782 = {1{`RANDOM}};
  windowBuffer_7 = _RAND_782[15:0];
  _RAND_783 = {1{`RANDOM}};
  windowBuffer_8 = _RAND_783[15:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      stateReg <= 2'h0;
    end else if (_T) begin
      if (io_enq_valid) begin
        stateReg <= 2'h1;
      end
    end else if (_T_1) begin
      if (_T_3) begin
        stateReg <= 2'h0;
      end else if (_T_4) begin
        stateReg <= 2'h1;
      end else if (_T_6) begin
        stateReg <= 2'h2;
      end
    end else if (_T_7) begin
      if (io_deq_ready) begin
        stateReg <= 2'h1;
      end
    end else if (_T_8) begin
      stateReg <= 2'h0;
    end
    if (_T) begin
      if (io_enq_valid) begin
        dataReg <= io_enq_bits;
      end
    end else if (_T_1) begin
      if (!(_T_3)) begin
        if (_T_4) begin
          dataReg <= io_enq_bits;
        end
      end
    end else if (_T_7) begin
      if (io_deq_ready) begin
        dataReg <= shadowReg;
      end
    end
    if (!(_T)) begin
      if (_T_1) begin
        if (!(_T_3)) begin
          if (!(_T_4)) begin
            if (_T_6) begin
              shadowReg <= io_enq_bits;
            end
          end
        end
      end
    end
    if (_T) begin
      userReg <= io_enq_user;
    end else if (_T_1) begin
      if (_T_3) begin
        userReg <= io_enq_user;
      end else if (_T_4) begin
        userReg <= io_enq_user;
      end
    end else if (_T_7) begin
      if (io_deq_ready) begin
        userReg <= shadowUserReg;
      end
    end
    if (!(_T)) begin
      if (_T_1) begin
        if (!(_T_3)) begin
          if (!(_T_4)) begin
            if (_T_6) begin
              shadowUserReg <= io_enq_user;
            end
          end
        end
      end
    end
    if (_T) begin
      if (io_enq_valid) begin
        lastReg <= io_enq_last;
      end
    end else if (_T_1) begin
      if (!(_T_3)) begin
        if (_T_4) begin
          lastReg <= io_enq_last;
        end
      end
    end else if (_T_7) begin
      if (io_deq_ready) begin
        lastReg <= shadowLastReg;
      end
    end
    if (!(_T)) begin
      if (_T_1) begin
        if (!(_T_3)) begin
          if (!(_T_4)) begin
            if (_T_6) begin
              shadowLastReg <= io_enq_last;
            end
          end
        end
      end
    end
    if (sel) begin
      lineBuffer_0 <= dataReg;
    end
    if (sel) begin
      lineBuffer_1 <= lineBuffer_0;
    end
    if (sel) begin
      lineBuffer_2 <= lineBuffer_1;
    end
    if (sel) begin
      lineBuffer_3 <= lineBuffer_2;
    end
    if (sel) begin
      lineBuffer_4 <= lineBuffer_3;
    end
    if (sel) begin
      lineBuffer_5 <= lineBuffer_4;
    end
    if (sel) begin
      lineBuffer_6 <= lineBuffer_5;
    end
    if (sel) begin
      lineBuffer_7 <= lineBuffer_6;
    end
    if (sel) begin
      lineBuffer_8 <= lineBuffer_7;
    end
    if (sel) begin
      lineBuffer_9 <= lineBuffer_8;
    end
    if (sel) begin
      lineBuffer_10 <= lineBuffer_9;
    end
    if (sel) begin
      lineBuffer_11 <= lineBuffer_10;
    end
    if (sel) begin
      lineBuffer_12 <= lineBuffer_11;
    end
    if (sel) begin
      lineBuffer_13 <= lineBuffer_12;
    end
    if (sel) begin
      lineBuffer_14 <= lineBuffer_13;
    end
    if (sel) begin
      lineBuffer_15 <= lineBuffer_14;
    end
    if (sel) begin
      lineBuffer_16 <= lineBuffer_15;
    end
    if (sel) begin
      lineBuffer_17 <= lineBuffer_16;
    end
    if (sel) begin
      lineBuffer_18 <= lineBuffer_17;
    end
    if (sel) begin
      lineBuffer_19 <= lineBuffer_18;
    end
    if (sel) begin
      lineBuffer_20 <= lineBuffer_19;
    end
    if (sel) begin
      lineBuffer_21 <= lineBuffer_20;
    end
    if (sel) begin
      lineBuffer_22 <= lineBuffer_21;
    end
    if (sel) begin
      lineBuffer_23 <= lineBuffer_22;
    end
    if (sel) begin
      lineBuffer_24 <= lineBuffer_23;
    end
    if (sel) begin
      lineBuffer_25 <= lineBuffer_24;
    end
    if (sel) begin
      lineBuffer_26 <= lineBuffer_25;
    end
    if (sel) begin
      lineBuffer_27 <= lineBuffer_26;
    end
    if (sel) begin
      lineBuffer_28 <= lineBuffer_27;
    end
    if (sel) begin
      lineBuffer_29 <= lineBuffer_28;
    end
    if (sel) begin
      lineBuffer_30 <= lineBuffer_29;
    end
    if (sel) begin
      lineBuffer_31 <= lineBuffer_30;
    end
    if (sel) begin
      lineBuffer_32 <= lineBuffer_31;
    end
    if (sel) begin
      lineBuffer_33 <= lineBuffer_32;
    end
    if (sel) begin
      lineBuffer_34 <= lineBuffer_33;
    end
    if (sel) begin
      lineBuffer_35 <= lineBuffer_34;
    end
    if (sel) begin
      lineBuffer_36 <= lineBuffer_35;
    end
    if (sel) begin
      lineBuffer_37 <= lineBuffer_36;
    end
    if (sel) begin
      lineBuffer_38 <= lineBuffer_37;
    end
    if (sel) begin
      lineBuffer_39 <= lineBuffer_38;
    end
    if (sel) begin
      lineBuffer_40 <= lineBuffer_39;
    end
    if (sel) begin
      lineBuffer_41 <= lineBuffer_40;
    end
    if (sel) begin
      lineBuffer_42 <= lineBuffer_41;
    end
    if (sel) begin
      lineBuffer_43 <= lineBuffer_42;
    end
    if (sel) begin
      lineBuffer_44 <= lineBuffer_43;
    end
    if (sel) begin
      lineBuffer_45 <= lineBuffer_44;
    end
    if (sel) begin
      lineBuffer_46 <= lineBuffer_45;
    end
    if (sel) begin
      lineBuffer_47 <= lineBuffer_46;
    end
    if (sel) begin
      lineBuffer_48 <= lineBuffer_47;
    end
    if (sel) begin
      lineBuffer_49 <= lineBuffer_48;
    end
    if (sel) begin
      lineBuffer_50 <= lineBuffer_49;
    end
    if (sel) begin
      lineBuffer_51 <= lineBuffer_50;
    end
    if (sel) begin
      lineBuffer_52 <= lineBuffer_51;
    end
    if (sel) begin
      lineBuffer_53 <= lineBuffer_52;
    end
    if (sel) begin
      lineBuffer_54 <= lineBuffer_53;
    end
    if (sel) begin
      lineBuffer_55 <= lineBuffer_54;
    end
    if (sel) begin
      lineBuffer_56 <= lineBuffer_55;
    end
    if (sel) begin
      lineBuffer_57 <= lineBuffer_56;
    end
    if (sel) begin
      lineBuffer_58 <= lineBuffer_57;
    end
    if (sel) begin
      lineBuffer_59 <= lineBuffer_58;
    end
    if (sel) begin
      lineBuffer_60 <= lineBuffer_59;
    end
    if (sel) begin
      lineBuffer_61 <= lineBuffer_60;
    end
    if (sel) begin
      lineBuffer_62 <= lineBuffer_61;
    end
    if (sel) begin
      lineBuffer_63 <= lineBuffer_62;
    end
    if (sel) begin
      lineBuffer_64 <= lineBuffer_63;
    end
    if (sel) begin
      lineBuffer_65 <= lineBuffer_64;
    end
    if (sel) begin
      lineBuffer_66 <= lineBuffer_65;
    end
    if (sel) begin
      lineBuffer_67 <= lineBuffer_66;
    end
    if (sel) begin
      lineBuffer_68 <= lineBuffer_67;
    end
    if (sel) begin
      lineBuffer_69 <= lineBuffer_68;
    end
    if (sel) begin
      lineBuffer_70 <= lineBuffer_69;
    end
    if (sel) begin
      lineBuffer_71 <= lineBuffer_70;
    end
    if (sel) begin
      lineBuffer_72 <= lineBuffer_71;
    end
    if (sel) begin
      lineBuffer_73 <= lineBuffer_72;
    end
    if (sel) begin
      lineBuffer_74 <= lineBuffer_73;
    end
    if (sel) begin
      lineBuffer_75 <= lineBuffer_74;
    end
    if (sel) begin
      lineBuffer_76 <= lineBuffer_75;
    end
    if (sel) begin
      lineBuffer_77 <= lineBuffer_76;
    end
    if (sel) begin
      lineBuffer_78 <= lineBuffer_77;
    end
    if (sel) begin
      lineBuffer_79 <= lineBuffer_78;
    end
    if (sel) begin
      lineBuffer_80 <= lineBuffer_79;
    end
    if (sel) begin
      lineBuffer_81 <= lineBuffer_80;
    end
    if (sel) begin
      lineBuffer_82 <= lineBuffer_81;
    end
    if (sel) begin
      lineBuffer_83 <= lineBuffer_82;
    end
    if (sel) begin
      lineBuffer_84 <= lineBuffer_83;
    end
    if (sel) begin
      lineBuffer_85 <= lineBuffer_84;
    end
    if (sel) begin
      lineBuffer_86 <= lineBuffer_85;
    end
    if (sel) begin
      lineBuffer_87 <= lineBuffer_86;
    end
    if (sel) begin
      lineBuffer_88 <= lineBuffer_87;
    end
    if (sel) begin
      lineBuffer_89 <= lineBuffer_88;
    end
    if (sel) begin
      lineBuffer_90 <= lineBuffer_89;
    end
    if (sel) begin
      lineBuffer_91 <= lineBuffer_90;
    end
    if (sel) begin
      lineBuffer_92 <= lineBuffer_91;
    end
    if (sel) begin
      lineBuffer_93 <= lineBuffer_92;
    end
    if (sel) begin
      lineBuffer_94 <= lineBuffer_93;
    end
    if (sel) begin
      lineBuffer_95 <= lineBuffer_94;
    end
    if (sel) begin
      lineBuffer_96 <= lineBuffer_95;
    end
    if (sel) begin
      lineBuffer_97 <= lineBuffer_96;
    end
    if (sel) begin
      lineBuffer_98 <= lineBuffer_97;
    end
    if (sel) begin
      lineBuffer_99 <= lineBuffer_98;
    end
    if (sel) begin
      lineBuffer_100 <= lineBuffer_99;
    end
    if (sel) begin
      lineBuffer_101 <= lineBuffer_100;
    end
    if (sel) begin
      lineBuffer_102 <= lineBuffer_101;
    end
    if (sel) begin
      lineBuffer_103 <= lineBuffer_102;
    end
    if (sel) begin
      lineBuffer_104 <= lineBuffer_103;
    end
    if (sel) begin
      lineBuffer_105 <= lineBuffer_104;
    end
    if (sel) begin
      lineBuffer_106 <= lineBuffer_105;
    end
    if (sel) begin
      lineBuffer_107 <= lineBuffer_106;
    end
    if (sel) begin
      lineBuffer_108 <= lineBuffer_107;
    end
    if (sel) begin
      lineBuffer_109 <= lineBuffer_108;
    end
    if (sel) begin
      lineBuffer_110 <= lineBuffer_109;
    end
    if (sel) begin
      lineBuffer_111 <= lineBuffer_110;
    end
    if (sel) begin
      lineBuffer_112 <= lineBuffer_111;
    end
    if (sel) begin
      lineBuffer_113 <= lineBuffer_112;
    end
    if (sel) begin
      lineBuffer_114 <= lineBuffer_113;
    end
    if (sel) begin
      lineBuffer_115 <= lineBuffer_114;
    end
    if (sel) begin
      lineBuffer_116 <= lineBuffer_115;
    end
    if (sel) begin
      lineBuffer_117 <= lineBuffer_116;
    end
    if (sel) begin
      lineBuffer_118 <= lineBuffer_117;
    end
    if (sel) begin
      lineBuffer_119 <= lineBuffer_118;
    end
    if (sel) begin
      lineBuffer_120 <= lineBuffer_119;
    end
    if (sel) begin
      lineBuffer_121 <= lineBuffer_120;
    end
    if (sel) begin
      lineBuffer_122 <= lineBuffer_121;
    end
    if (sel) begin
      lineBuffer_123 <= lineBuffer_122;
    end
    if (sel) begin
      lineBuffer_124 <= lineBuffer_123;
    end
    if (sel) begin
      lineBuffer_125 <= lineBuffer_124;
    end
    if (sel) begin
      lineBuffer_126 <= lineBuffer_125;
    end
    if (sel) begin
      lineBuffer_127 <= lineBuffer_126;
    end
    if (sel) begin
      lineBuffer_128 <= lineBuffer_127;
    end
    if (sel) begin
      lineBuffer_129 <= lineBuffer_128;
    end
    if (sel) begin
      lineBuffer_130 <= lineBuffer_129;
    end
    if (sel) begin
      lineBuffer_131 <= lineBuffer_130;
    end
    if (sel) begin
      lineBuffer_132 <= lineBuffer_131;
    end
    if (sel) begin
      lineBuffer_133 <= lineBuffer_132;
    end
    if (sel) begin
      lineBuffer_134 <= lineBuffer_133;
    end
    if (sel) begin
      lineBuffer_135 <= lineBuffer_134;
    end
    if (sel) begin
      lineBuffer_136 <= lineBuffer_135;
    end
    if (sel) begin
      lineBuffer_137 <= lineBuffer_136;
    end
    if (sel) begin
      lineBuffer_138 <= lineBuffer_137;
    end
    if (sel) begin
      lineBuffer_139 <= lineBuffer_138;
    end
    if (sel) begin
      lineBuffer_140 <= lineBuffer_139;
    end
    if (sel) begin
      lineBuffer_141 <= lineBuffer_140;
    end
    if (sel) begin
      lineBuffer_142 <= lineBuffer_141;
    end
    if (sel) begin
      lineBuffer_143 <= lineBuffer_142;
    end
    if (sel) begin
      lineBuffer_144 <= lineBuffer_143;
    end
    if (sel) begin
      lineBuffer_145 <= lineBuffer_144;
    end
    if (sel) begin
      lineBuffer_146 <= lineBuffer_145;
    end
    if (sel) begin
      lineBuffer_147 <= lineBuffer_146;
    end
    if (sel) begin
      lineBuffer_148 <= lineBuffer_147;
    end
    if (sel) begin
      lineBuffer_149 <= lineBuffer_148;
    end
    if (sel) begin
      lineBuffer_150 <= lineBuffer_149;
    end
    if (sel) begin
      lineBuffer_151 <= lineBuffer_150;
    end
    if (sel) begin
      lineBuffer_152 <= lineBuffer_151;
    end
    if (sel) begin
      lineBuffer_153 <= lineBuffer_152;
    end
    if (sel) begin
      lineBuffer_154 <= lineBuffer_153;
    end
    if (sel) begin
      lineBuffer_155 <= lineBuffer_154;
    end
    if (sel) begin
      lineBuffer_156 <= lineBuffer_155;
    end
    if (sel) begin
      lineBuffer_157 <= lineBuffer_156;
    end
    if (sel) begin
      lineBuffer_158 <= lineBuffer_157;
    end
    if (sel) begin
      lineBuffer_159 <= lineBuffer_158;
    end
    if (sel) begin
      lineBuffer_160 <= lineBuffer_159;
    end
    if (sel) begin
      lineBuffer_161 <= lineBuffer_160;
    end
    if (sel) begin
      lineBuffer_162 <= lineBuffer_161;
    end
    if (sel) begin
      lineBuffer_163 <= lineBuffer_162;
    end
    if (sel) begin
      lineBuffer_164 <= lineBuffer_163;
    end
    if (sel) begin
      lineBuffer_165 <= lineBuffer_164;
    end
    if (sel) begin
      lineBuffer_166 <= lineBuffer_165;
    end
    if (sel) begin
      lineBuffer_167 <= lineBuffer_166;
    end
    if (sel) begin
      lineBuffer_168 <= lineBuffer_167;
    end
    if (sel) begin
      lineBuffer_169 <= lineBuffer_168;
    end
    if (sel) begin
      lineBuffer_170 <= lineBuffer_169;
    end
    if (sel) begin
      lineBuffer_171 <= lineBuffer_170;
    end
    if (sel) begin
      lineBuffer_172 <= lineBuffer_171;
    end
    if (sel) begin
      lineBuffer_173 <= lineBuffer_172;
    end
    if (sel) begin
      lineBuffer_174 <= lineBuffer_173;
    end
    if (sel) begin
      lineBuffer_175 <= lineBuffer_174;
    end
    if (sel) begin
      lineBuffer_176 <= lineBuffer_175;
    end
    if (sel) begin
      lineBuffer_177 <= lineBuffer_176;
    end
    if (sel) begin
      lineBuffer_178 <= lineBuffer_177;
    end
    if (sel) begin
      lineBuffer_179 <= lineBuffer_178;
    end
    if (sel) begin
      lineBuffer_180 <= lineBuffer_179;
    end
    if (sel) begin
      lineBuffer_181 <= lineBuffer_180;
    end
    if (sel) begin
      lineBuffer_182 <= lineBuffer_181;
    end
    if (sel) begin
      lineBuffer_183 <= lineBuffer_182;
    end
    if (sel) begin
      lineBuffer_184 <= lineBuffer_183;
    end
    if (sel) begin
      lineBuffer_185 <= lineBuffer_184;
    end
    if (sel) begin
      lineBuffer_186 <= lineBuffer_185;
    end
    if (sel) begin
      lineBuffer_187 <= lineBuffer_186;
    end
    if (sel) begin
      lineBuffer_188 <= lineBuffer_187;
    end
    if (sel) begin
      lineBuffer_189 <= lineBuffer_188;
    end
    if (sel) begin
      lineBuffer_190 <= lineBuffer_189;
    end
    if (sel) begin
      lineBuffer_191 <= lineBuffer_190;
    end
    if (sel) begin
      lineBuffer_192 <= lineBuffer_191;
    end
    if (sel) begin
      lineBuffer_193 <= lineBuffer_192;
    end
    if (sel) begin
      lineBuffer_194 <= lineBuffer_193;
    end
    if (sel) begin
      lineBuffer_195 <= lineBuffer_194;
    end
    if (sel) begin
      lineBuffer_196 <= lineBuffer_195;
    end
    if (sel) begin
      lineBuffer_197 <= lineBuffer_196;
    end
    if (sel) begin
      lineBuffer_198 <= lineBuffer_197;
    end
    if (sel) begin
      lineBuffer_199 <= lineBuffer_198;
    end
    if (sel) begin
      lineBuffer_200 <= lineBuffer_199;
    end
    if (sel) begin
      lineBuffer_201 <= lineBuffer_200;
    end
    if (sel) begin
      lineBuffer_202 <= lineBuffer_201;
    end
    if (sel) begin
      lineBuffer_203 <= lineBuffer_202;
    end
    if (sel) begin
      lineBuffer_204 <= lineBuffer_203;
    end
    if (sel) begin
      lineBuffer_205 <= lineBuffer_204;
    end
    if (sel) begin
      lineBuffer_206 <= lineBuffer_205;
    end
    if (sel) begin
      lineBuffer_207 <= lineBuffer_206;
    end
    if (sel) begin
      lineBuffer_208 <= lineBuffer_207;
    end
    if (sel) begin
      lineBuffer_209 <= lineBuffer_208;
    end
    if (sel) begin
      lineBuffer_210 <= lineBuffer_209;
    end
    if (sel) begin
      lineBuffer_211 <= lineBuffer_210;
    end
    if (sel) begin
      lineBuffer_212 <= lineBuffer_211;
    end
    if (sel) begin
      lineBuffer_213 <= lineBuffer_212;
    end
    if (sel) begin
      lineBuffer_214 <= lineBuffer_213;
    end
    if (sel) begin
      lineBuffer_215 <= lineBuffer_214;
    end
    if (sel) begin
      lineBuffer_216 <= lineBuffer_215;
    end
    if (sel) begin
      lineBuffer_217 <= lineBuffer_216;
    end
    if (sel) begin
      lineBuffer_218 <= lineBuffer_217;
    end
    if (sel) begin
      lineBuffer_219 <= lineBuffer_218;
    end
    if (sel) begin
      lineBuffer_220 <= lineBuffer_219;
    end
    if (sel) begin
      lineBuffer_221 <= lineBuffer_220;
    end
    if (sel) begin
      lineBuffer_222 <= lineBuffer_221;
    end
    if (sel) begin
      lineBuffer_223 <= lineBuffer_222;
    end
    if (sel) begin
      lineBuffer_224 <= lineBuffer_223;
    end
    if (sel) begin
      lineBuffer_225 <= lineBuffer_224;
    end
    if (sel) begin
      lineBuffer_226 <= lineBuffer_225;
    end
    if (sel) begin
      lineBuffer_227 <= lineBuffer_226;
    end
    if (sel) begin
      lineBuffer_228 <= lineBuffer_227;
    end
    if (sel) begin
      lineBuffer_229 <= lineBuffer_228;
    end
    if (sel) begin
      lineBuffer_230 <= lineBuffer_229;
    end
    if (sel) begin
      lineBuffer_231 <= lineBuffer_230;
    end
    if (sel) begin
      lineBuffer_232 <= lineBuffer_231;
    end
    if (sel) begin
      lineBuffer_233 <= lineBuffer_232;
    end
    if (sel) begin
      lineBuffer_234 <= lineBuffer_233;
    end
    if (sel) begin
      lineBuffer_235 <= lineBuffer_234;
    end
    if (sel) begin
      lineBuffer_236 <= lineBuffer_235;
    end
    if (sel) begin
      lineBuffer_237 <= lineBuffer_236;
    end
    if (sel) begin
      lineBuffer_238 <= lineBuffer_237;
    end
    if (sel) begin
      lineBuffer_239 <= lineBuffer_238;
    end
    if (sel) begin
      lineBuffer_240 <= lineBuffer_239;
    end
    if (sel) begin
      lineBuffer_241 <= lineBuffer_240;
    end
    if (sel) begin
      lineBuffer_242 <= lineBuffer_241;
    end
    if (sel) begin
      lineBuffer_243 <= lineBuffer_242;
    end
    if (sel) begin
      lineBuffer_244 <= lineBuffer_243;
    end
    if (sel) begin
      lineBuffer_245 <= lineBuffer_244;
    end
    if (sel) begin
      lineBuffer_246 <= lineBuffer_245;
    end
    if (sel) begin
      lineBuffer_247 <= lineBuffer_246;
    end
    if (sel) begin
      lineBuffer_248 <= lineBuffer_247;
    end
    if (sel) begin
      lineBuffer_249 <= lineBuffer_248;
    end
    if (sel) begin
      lineBuffer_250 <= lineBuffer_249;
    end
    if (sel) begin
      lineBuffer_251 <= lineBuffer_250;
    end
    if (sel) begin
      lineBuffer_252 <= lineBuffer_251;
    end
    if (sel) begin
      lineBuffer_253 <= lineBuffer_252;
    end
    if (sel) begin
      lineBuffer_254 <= lineBuffer_253;
    end
    if (sel) begin
      lineBuffer_255 <= lineBuffer_254;
    end
    if (sel) begin
      lineBuffer_256 <= lineBuffer_255;
    end
    if (sel) begin
      lineBuffer_257 <= lineBuffer_256;
    end
    if (sel) begin
      lineBuffer_258 <= lineBuffer_257;
    end
    if (sel) begin
      lineBuffer_259 <= lineBuffer_258;
    end
    if (sel) begin
      lineBuffer_260 <= lineBuffer_259;
    end
    if (sel) begin
      lineBuffer_261 <= lineBuffer_260;
    end
    if (sel) begin
      lineBuffer_262 <= lineBuffer_261;
    end
    if (sel) begin
      lineBuffer_263 <= lineBuffer_262;
    end
    if (sel) begin
      lineBuffer_264 <= lineBuffer_263;
    end
    if (sel) begin
      lineBuffer_265 <= lineBuffer_264;
    end
    if (sel) begin
      lineBuffer_266 <= lineBuffer_265;
    end
    if (sel) begin
      lineBuffer_267 <= lineBuffer_266;
    end
    if (sel) begin
      lineBuffer_268 <= lineBuffer_267;
    end
    if (sel) begin
      lineBuffer_269 <= lineBuffer_268;
    end
    if (sel) begin
      lineBuffer_270 <= lineBuffer_269;
    end
    if (sel) begin
      lineBuffer_271 <= lineBuffer_270;
    end
    if (sel) begin
      lineBuffer_272 <= lineBuffer_271;
    end
    if (sel) begin
      lineBuffer_273 <= lineBuffer_272;
    end
    if (sel) begin
      lineBuffer_274 <= lineBuffer_273;
    end
    if (sel) begin
      lineBuffer_275 <= lineBuffer_274;
    end
    if (sel) begin
      lineBuffer_276 <= lineBuffer_275;
    end
    if (sel) begin
      lineBuffer_277 <= lineBuffer_276;
    end
    if (sel) begin
      lineBuffer_278 <= lineBuffer_277;
    end
    if (sel) begin
      lineBuffer_279 <= lineBuffer_278;
    end
    if (sel) begin
      lineBuffer_280 <= lineBuffer_279;
    end
    if (sel) begin
      lineBuffer_281 <= lineBuffer_280;
    end
    if (sel) begin
      lineBuffer_282 <= lineBuffer_281;
    end
    if (sel) begin
      lineBuffer_283 <= lineBuffer_282;
    end
    if (sel) begin
      lineBuffer_284 <= lineBuffer_283;
    end
    if (sel) begin
      lineBuffer_285 <= lineBuffer_284;
    end
    if (sel) begin
      lineBuffer_286 <= lineBuffer_285;
    end
    if (sel) begin
      lineBuffer_287 <= lineBuffer_286;
    end
    if (sel) begin
      lineBuffer_288 <= lineBuffer_287;
    end
    if (sel) begin
      lineBuffer_289 <= lineBuffer_288;
    end
    if (sel) begin
      lineBuffer_290 <= lineBuffer_289;
    end
    if (sel) begin
      lineBuffer_291 <= lineBuffer_290;
    end
    if (sel) begin
      lineBuffer_292 <= lineBuffer_291;
    end
    if (sel) begin
      lineBuffer_293 <= lineBuffer_292;
    end
    if (sel) begin
      lineBuffer_294 <= lineBuffer_293;
    end
    if (sel) begin
      lineBuffer_295 <= lineBuffer_294;
    end
    if (sel) begin
      lineBuffer_296 <= lineBuffer_295;
    end
    if (sel) begin
      lineBuffer_297 <= lineBuffer_296;
    end
    if (sel) begin
      lineBuffer_298 <= lineBuffer_297;
    end
    if (sel) begin
      lineBuffer_299 <= lineBuffer_298;
    end
    if (sel) begin
      lineBuffer_300 <= lineBuffer_299;
    end
    if (sel) begin
      lineBuffer_301 <= lineBuffer_300;
    end
    if (sel) begin
      lineBuffer_302 <= lineBuffer_301;
    end
    if (sel) begin
      lineBuffer_303 <= lineBuffer_302;
    end
    if (sel) begin
      lineBuffer_304 <= lineBuffer_303;
    end
    if (sel) begin
      lineBuffer_305 <= lineBuffer_304;
    end
    if (sel) begin
      lineBuffer_306 <= lineBuffer_305;
    end
    if (sel) begin
      lineBuffer_307 <= lineBuffer_306;
    end
    if (sel) begin
      lineBuffer_308 <= lineBuffer_307;
    end
    if (sel) begin
      lineBuffer_309 <= lineBuffer_308;
    end
    if (sel) begin
      lineBuffer_310 <= lineBuffer_309;
    end
    if (sel) begin
      lineBuffer_311 <= lineBuffer_310;
    end
    if (sel) begin
      lineBuffer_312 <= lineBuffer_311;
    end
    if (sel) begin
      lineBuffer_313 <= lineBuffer_312;
    end
    if (sel) begin
      lineBuffer_314 <= lineBuffer_313;
    end
    if (sel) begin
      lineBuffer_315 <= lineBuffer_314;
    end
    if (sel) begin
      lineBuffer_316 <= lineBuffer_315;
    end
    if (sel) begin
      lineBuffer_317 <= lineBuffer_316;
    end
    if (sel) begin
      lineBuffer_318 <= lineBuffer_317;
    end
    if (sel) begin
      lineBuffer_319 <= lineBuffer_318;
    end
    if (sel) begin
      lineBuffer_320 <= lineBuffer_319;
    end
    if (sel) begin
      lineBuffer_321 <= lineBuffer_320;
    end
    if (sel) begin
      lineBuffer_322 <= lineBuffer_321;
    end
    if (sel) begin
      lineBuffer_323 <= lineBuffer_322;
    end
    if (sel) begin
      lineBuffer_324 <= lineBuffer_323;
    end
    if (sel) begin
      lineBuffer_325 <= lineBuffer_324;
    end
    if (sel) begin
      lineBuffer_326 <= lineBuffer_325;
    end
    if (sel) begin
      lineBuffer_327 <= lineBuffer_326;
    end
    if (sel) begin
      lineBuffer_328 <= lineBuffer_327;
    end
    if (sel) begin
      lineBuffer_329 <= lineBuffer_328;
    end
    if (sel) begin
      lineBuffer_330 <= lineBuffer_329;
    end
    if (sel) begin
      lineBuffer_331 <= lineBuffer_330;
    end
    if (sel) begin
      lineBuffer_332 <= lineBuffer_331;
    end
    if (sel) begin
      lineBuffer_333 <= lineBuffer_332;
    end
    if (sel) begin
      lineBuffer_334 <= lineBuffer_333;
    end
    if (sel) begin
      lineBuffer_335 <= lineBuffer_334;
    end
    if (sel) begin
      lineBuffer_336 <= lineBuffer_335;
    end
    if (sel) begin
      lineBuffer_337 <= lineBuffer_336;
    end
    if (sel) begin
      lineBuffer_338 <= lineBuffer_337;
    end
    if (sel) begin
      lineBuffer_339 <= lineBuffer_338;
    end
    if (sel) begin
      lineBuffer_340 <= lineBuffer_339;
    end
    if (sel) begin
      lineBuffer_341 <= lineBuffer_340;
    end
    if (sel) begin
      lineBuffer_342 <= lineBuffer_341;
    end
    if (sel) begin
      lineBuffer_343 <= lineBuffer_342;
    end
    if (sel) begin
      lineBuffer_344 <= lineBuffer_343;
    end
    if (sel) begin
      lineBuffer_345 <= lineBuffer_344;
    end
    if (sel) begin
      lineBuffer_346 <= lineBuffer_345;
    end
    if (sel) begin
      lineBuffer_347 <= lineBuffer_346;
    end
    if (sel) begin
      lineBuffer_348 <= lineBuffer_347;
    end
    if (sel) begin
      lineBuffer_349 <= lineBuffer_348;
    end
    if (sel) begin
      lineBuffer_350 <= lineBuffer_349;
    end
    if (sel) begin
      lineBuffer_351 <= lineBuffer_350;
    end
    if (sel) begin
      lineBuffer_352 <= lineBuffer_351;
    end
    if (sel) begin
      lineBuffer_353 <= lineBuffer_352;
    end
    if (sel) begin
      lineBuffer_354 <= lineBuffer_353;
    end
    if (sel) begin
      lineBuffer_355 <= lineBuffer_354;
    end
    if (sel) begin
      lineBuffer_356 <= lineBuffer_355;
    end
    if (sel) begin
      lineBuffer_357 <= lineBuffer_356;
    end
    if (sel) begin
      lineBuffer_358 <= lineBuffer_357;
    end
    if (sel) begin
      lineBuffer_359 <= lineBuffer_358;
    end
    if (sel) begin
      lineBuffer_360 <= lineBuffer_359;
    end
    if (sel) begin
      lineBuffer_361 <= lineBuffer_360;
    end
    if (sel) begin
      lineBuffer_362 <= lineBuffer_361;
    end
    if (sel) begin
      lineBuffer_363 <= lineBuffer_362;
    end
    if (sel) begin
      lineBuffer_364 <= lineBuffer_363;
    end
    if (sel) begin
      lineBuffer_365 <= lineBuffer_364;
    end
    if (sel) begin
      lineBuffer_366 <= lineBuffer_365;
    end
    if (sel) begin
      lineBuffer_367 <= lineBuffer_366;
    end
    if (sel) begin
      lineBuffer_368 <= lineBuffer_367;
    end
    if (sel) begin
      lineBuffer_369 <= lineBuffer_368;
    end
    if (sel) begin
      lineBuffer_370 <= lineBuffer_369;
    end
    if (sel) begin
      lineBuffer_371 <= lineBuffer_370;
    end
    if (sel) begin
      lineBuffer_372 <= lineBuffer_371;
    end
    if (sel) begin
      lineBuffer_373 <= lineBuffer_372;
    end
    if (sel) begin
      lineBuffer_374 <= lineBuffer_373;
    end
    if (sel) begin
      lineBuffer_375 <= lineBuffer_374;
    end
    if (sel) begin
      lineBuffer_376 <= lineBuffer_375;
    end
    if (sel) begin
      lineBuffer_377 <= lineBuffer_376;
    end
    if (sel) begin
      lineBuffer_378 <= lineBuffer_377;
    end
    if (sel) begin
      lineBuffer_379 <= lineBuffer_378;
    end
    if (sel) begin
      lineBuffer_380 <= lineBuffer_379;
    end
    if (sel) begin
      lineBuffer_381 <= lineBuffer_380;
    end
    if (sel) begin
      lineBuffer_382 <= lineBuffer_381;
    end
    if (sel) begin
      lineBuffer_383 <= lineBuffer_382;
    end
    if (sel) begin
      lineBuffer_384 <= lineBuffer_383;
    end
    if (sel) begin
      lineBuffer_385 <= lineBuffer_384;
    end
    if (sel) begin
      lineBuffer_386 <= lineBuffer_385;
    end
    if (sel) begin
      lineBuffer_387 <= lineBuffer_386;
    end
    if (sel) begin
      lineBuffer_388 <= lineBuffer_387;
    end
    if (sel) begin
      lineBuffer_389 <= lineBuffer_388;
    end
    if (sel) begin
      lineBuffer_390 <= lineBuffer_389;
    end
    if (sel) begin
      lineBuffer_391 <= lineBuffer_390;
    end
    if (sel) begin
      lineBuffer_392 <= lineBuffer_391;
    end
    if (sel) begin
      lineBuffer_393 <= lineBuffer_392;
    end
    if (sel) begin
      lineBuffer_394 <= lineBuffer_393;
    end
    if (sel) begin
      lineBuffer_395 <= lineBuffer_394;
    end
    if (sel) begin
      lineBuffer_396 <= lineBuffer_395;
    end
    if (sel) begin
      lineBuffer_397 <= lineBuffer_396;
    end
    if (sel) begin
      lineBuffer_398 <= lineBuffer_397;
    end
    if (sel) begin
      lineBuffer_399 <= lineBuffer_398;
    end
    if (sel) begin
      lineBuffer_400 <= lineBuffer_399;
    end
    if (sel) begin
      lineBuffer_401 <= lineBuffer_400;
    end
    if (sel) begin
      lineBuffer_402 <= lineBuffer_401;
    end
    if (sel) begin
      lineBuffer_403 <= lineBuffer_402;
    end
    if (sel) begin
      lineBuffer_404 <= lineBuffer_403;
    end
    if (sel) begin
      lineBuffer_405 <= lineBuffer_404;
    end
    if (sel) begin
      lineBuffer_406 <= lineBuffer_405;
    end
    if (sel) begin
      lineBuffer_407 <= lineBuffer_406;
    end
    if (sel) begin
      lineBuffer_408 <= lineBuffer_407;
    end
    if (sel) begin
      lineBuffer_409 <= lineBuffer_408;
    end
    if (sel) begin
      lineBuffer_410 <= lineBuffer_409;
    end
    if (sel) begin
      lineBuffer_411 <= lineBuffer_410;
    end
    if (sel) begin
      lineBuffer_412 <= lineBuffer_411;
    end
    if (sel) begin
      lineBuffer_413 <= lineBuffer_412;
    end
    if (sel) begin
      lineBuffer_414 <= lineBuffer_413;
    end
    if (sel) begin
      lineBuffer_415 <= lineBuffer_414;
    end
    if (sel) begin
      lineBuffer_416 <= lineBuffer_415;
    end
    if (sel) begin
      lineBuffer_417 <= lineBuffer_416;
    end
    if (sel) begin
      lineBuffer_418 <= lineBuffer_417;
    end
    if (sel) begin
      lineBuffer_419 <= lineBuffer_418;
    end
    if (sel) begin
      lineBuffer_420 <= lineBuffer_419;
    end
    if (sel) begin
      lineBuffer_421 <= lineBuffer_420;
    end
    if (sel) begin
      lineBuffer_422 <= lineBuffer_421;
    end
    if (sel) begin
      lineBuffer_423 <= lineBuffer_422;
    end
    if (sel) begin
      lineBuffer_424 <= lineBuffer_423;
    end
    if (sel) begin
      lineBuffer_425 <= lineBuffer_424;
    end
    if (sel) begin
      lineBuffer_426 <= lineBuffer_425;
    end
    if (sel) begin
      lineBuffer_427 <= lineBuffer_426;
    end
    if (sel) begin
      lineBuffer_428 <= lineBuffer_427;
    end
    if (sel) begin
      lineBuffer_429 <= lineBuffer_428;
    end
    if (sel) begin
      lineBuffer_430 <= lineBuffer_429;
    end
    if (sel) begin
      lineBuffer_431 <= lineBuffer_430;
    end
    if (sel) begin
      lineBuffer_432 <= lineBuffer_431;
    end
    if (sel) begin
      lineBuffer_433 <= lineBuffer_432;
    end
    if (sel) begin
      lineBuffer_434 <= lineBuffer_433;
    end
    if (sel) begin
      lineBuffer_435 <= lineBuffer_434;
    end
    if (sel) begin
      lineBuffer_436 <= lineBuffer_435;
    end
    if (sel) begin
      lineBuffer_437 <= lineBuffer_436;
    end
    if (sel) begin
      lineBuffer_438 <= lineBuffer_437;
    end
    if (sel) begin
      lineBuffer_439 <= lineBuffer_438;
    end
    if (sel) begin
      lineBuffer_440 <= lineBuffer_439;
    end
    if (sel) begin
      lineBuffer_441 <= lineBuffer_440;
    end
    if (sel) begin
      lineBuffer_442 <= lineBuffer_441;
    end
    if (sel) begin
      lineBuffer_443 <= lineBuffer_442;
    end
    if (sel) begin
      lineBuffer_444 <= lineBuffer_443;
    end
    if (sel) begin
      lineBuffer_445 <= lineBuffer_444;
    end
    if (sel) begin
      lineBuffer_446 <= lineBuffer_445;
    end
    if (sel) begin
      lineBuffer_447 <= lineBuffer_446;
    end
    if (sel) begin
      lineBuffer_448 <= lineBuffer_447;
    end
    if (sel) begin
      lineBuffer_449 <= lineBuffer_448;
    end
    if (sel) begin
      lineBuffer_450 <= lineBuffer_449;
    end
    if (sel) begin
      lineBuffer_451 <= lineBuffer_450;
    end
    if (sel) begin
      lineBuffer_452 <= lineBuffer_451;
    end
    if (sel) begin
      lineBuffer_453 <= lineBuffer_452;
    end
    if (sel) begin
      lineBuffer_454 <= lineBuffer_453;
    end
    if (sel) begin
      lineBuffer_455 <= lineBuffer_454;
    end
    if (sel) begin
      lineBuffer_456 <= lineBuffer_455;
    end
    if (sel) begin
      lineBuffer_457 <= lineBuffer_456;
    end
    if (sel) begin
      lineBuffer_458 <= lineBuffer_457;
    end
    if (sel) begin
      lineBuffer_459 <= lineBuffer_458;
    end
    if (sel) begin
      lineBuffer_460 <= lineBuffer_459;
    end
    if (sel) begin
      lineBuffer_461 <= lineBuffer_460;
    end
    if (sel) begin
      lineBuffer_462 <= lineBuffer_461;
    end
    if (sel) begin
      lineBuffer_463 <= lineBuffer_462;
    end
    if (sel) begin
      lineBuffer_464 <= lineBuffer_463;
    end
    if (sel) begin
      lineBuffer_465 <= lineBuffer_464;
    end
    if (sel) begin
      lineBuffer_466 <= lineBuffer_465;
    end
    if (sel) begin
      lineBuffer_467 <= lineBuffer_466;
    end
    if (sel) begin
      lineBuffer_468 <= lineBuffer_467;
    end
    if (sel) begin
      lineBuffer_469 <= lineBuffer_468;
    end
    if (sel) begin
      lineBuffer_470 <= lineBuffer_469;
    end
    if (sel) begin
      lineBuffer_471 <= lineBuffer_470;
    end
    if (sel) begin
      lineBuffer_472 <= lineBuffer_471;
    end
    if (sel) begin
      lineBuffer_473 <= lineBuffer_472;
    end
    if (sel) begin
      lineBuffer_474 <= lineBuffer_473;
    end
    if (sel) begin
      lineBuffer_475 <= lineBuffer_474;
    end
    if (sel) begin
      lineBuffer_476 <= lineBuffer_475;
    end
    if (sel) begin
      lineBuffer_477 <= lineBuffer_476;
    end
    if (sel) begin
      lineBuffer_478 <= lineBuffer_477;
    end
    if (sel) begin
      lineBuffer_479 <= lineBuffer_478;
    end
    if (sel) begin
      lineBuffer_480 <= lineBuffer_479;
    end
    if (sel) begin
      lineBuffer_481 <= lineBuffer_480;
    end
    if (sel) begin
      lineBuffer_482 <= lineBuffer_481;
    end
    if (sel) begin
      lineBuffer_483 <= lineBuffer_482;
    end
    if (sel) begin
      lineBuffer_484 <= lineBuffer_483;
    end
    if (sel) begin
      lineBuffer_485 <= lineBuffer_484;
    end
    if (sel) begin
      lineBuffer_486 <= lineBuffer_485;
    end
    if (sel) begin
      lineBuffer_487 <= lineBuffer_486;
    end
    if (sel) begin
      lineBuffer_488 <= lineBuffer_487;
    end
    if (sel) begin
      lineBuffer_489 <= lineBuffer_488;
    end
    if (sel) begin
      lineBuffer_490 <= lineBuffer_489;
    end
    if (sel) begin
      lineBuffer_491 <= lineBuffer_490;
    end
    if (sel) begin
      lineBuffer_492 <= lineBuffer_491;
    end
    if (sel) begin
      lineBuffer_493 <= lineBuffer_492;
    end
    if (sel) begin
      lineBuffer_494 <= lineBuffer_493;
    end
    if (sel) begin
      lineBuffer_495 <= lineBuffer_494;
    end
    if (sel) begin
      lineBuffer_496 <= lineBuffer_495;
    end
    if (sel) begin
      lineBuffer_497 <= lineBuffer_496;
    end
    if (sel) begin
      lineBuffer_498 <= lineBuffer_497;
    end
    if (sel) begin
      lineBuffer_499 <= lineBuffer_498;
    end
    if (sel) begin
      lineBuffer_500 <= lineBuffer_499;
    end
    if (sel) begin
      lineBuffer_501 <= lineBuffer_500;
    end
    if (sel) begin
      lineBuffer_502 <= lineBuffer_501;
    end
    if (sel) begin
      lineBuffer_503 <= lineBuffer_502;
    end
    if (sel) begin
      lineBuffer_504 <= lineBuffer_503;
    end
    if (sel) begin
      lineBuffer_505 <= lineBuffer_504;
    end
    if (sel) begin
      lineBuffer_506 <= lineBuffer_505;
    end
    if (sel) begin
      lineBuffer_507 <= lineBuffer_506;
    end
    if (sel) begin
      lineBuffer_508 <= lineBuffer_507;
    end
    if (sel) begin
      lineBuffer_509 <= lineBuffer_508;
    end
    if (sel) begin
      lineBuffer_510 <= lineBuffer_509;
    end
    if (sel) begin
      lineBuffer_511 <= lineBuffer_510;
    end
    if (sel) begin
      lineBuffer_512 <= lineBuffer_511;
    end
    if (sel) begin
      lineBuffer_513 <= lineBuffer_512;
    end
    if (sel) begin
      lineBuffer_514 <= lineBuffer_513;
    end
    if (sel) begin
      lineBuffer_515 <= lineBuffer_514;
    end
    if (sel) begin
      lineBuffer_516 <= lineBuffer_515;
    end
    if (sel) begin
      lineBuffer_517 <= lineBuffer_516;
    end
    if (sel) begin
      lineBuffer_518 <= lineBuffer_517;
    end
    if (sel) begin
      lineBuffer_519 <= lineBuffer_518;
    end
    if (sel) begin
      lineBuffer_520 <= lineBuffer_519;
    end
    if (sel) begin
      lineBuffer_521 <= lineBuffer_520;
    end
    if (sel) begin
      lineBuffer_522 <= lineBuffer_521;
    end
    if (sel) begin
      lineBuffer_523 <= lineBuffer_522;
    end
    if (sel) begin
      lineBuffer_524 <= lineBuffer_523;
    end
    if (sel) begin
      lineBuffer_525 <= lineBuffer_524;
    end
    if (sel) begin
      lineBuffer_526 <= lineBuffer_525;
    end
    if (sel) begin
      lineBuffer_527 <= lineBuffer_526;
    end
    if (sel) begin
      lineBuffer_528 <= lineBuffer_527;
    end
    if (sel) begin
      lineBuffer_529 <= lineBuffer_528;
    end
    if (sel) begin
      lineBuffer_530 <= lineBuffer_529;
    end
    if (sel) begin
      lineBuffer_531 <= lineBuffer_530;
    end
    if (sel) begin
      lineBuffer_532 <= lineBuffer_531;
    end
    if (sel) begin
      lineBuffer_533 <= lineBuffer_532;
    end
    if (sel) begin
      lineBuffer_534 <= lineBuffer_533;
    end
    if (sel) begin
      lineBuffer_535 <= lineBuffer_534;
    end
    if (sel) begin
      lineBuffer_536 <= lineBuffer_535;
    end
    if (sel) begin
      lineBuffer_537 <= lineBuffer_536;
    end
    if (sel) begin
      lineBuffer_538 <= lineBuffer_537;
    end
    if (sel) begin
      lineBuffer_539 <= lineBuffer_538;
    end
    if (sel) begin
      lineBuffer_540 <= lineBuffer_539;
    end
    if (sel) begin
      lineBuffer_541 <= lineBuffer_540;
    end
    if (sel) begin
      lineBuffer_542 <= lineBuffer_541;
    end
    if (sel) begin
      lineBuffer_543 <= lineBuffer_542;
    end
    if (sel) begin
      lineBuffer_544 <= lineBuffer_543;
    end
    if (sel) begin
      lineBuffer_545 <= lineBuffer_544;
    end
    if (sel) begin
      lineBuffer_546 <= lineBuffer_545;
    end
    if (sel) begin
      lineBuffer_547 <= lineBuffer_546;
    end
    if (sel) begin
      lineBuffer_548 <= lineBuffer_547;
    end
    if (sel) begin
      lineBuffer_549 <= lineBuffer_548;
    end
    if (sel) begin
      lineBuffer_550 <= lineBuffer_549;
    end
    if (sel) begin
      lineBuffer_551 <= lineBuffer_550;
    end
    if (sel) begin
      lineBuffer_552 <= lineBuffer_551;
    end
    if (sel) begin
      lineBuffer_553 <= lineBuffer_552;
    end
    if (sel) begin
      lineBuffer_554 <= lineBuffer_553;
    end
    if (sel) begin
      lineBuffer_555 <= lineBuffer_554;
    end
    if (sel) begin
      lineBuffer_556 <= lineBuffer_555;
    end
    if (sel) begin
      lineBuffer_557 <= lineBuffer_556;
    end
    if (sel) begin
      lineBuffer_558 <= lineBuffer_557;
    end
    if (sel) begin
      lineBuffer_559 <= lineBuffer_558;
    end
    if (sel) begin
      lineBuffer_560 <= lineBuffer_559;
    end
    if (sel) begin
      lineBuffer_561 <= lineBuffer_560;
    end
    if (sel) begin
      lineBuffer_562 <= lineBuffer_561;
    end
    if (sel) begin
      lineBuffer_563 <= lineBuffer_562;
    end
    if (sel) begin
      lineBuffer_564 <= lineBuffer_563;
    end
    if (sel) begin
      lineBuffer_565 <= lineBuffer_564;
    end
    if (sel) begin
      lineBuffer_566 <= lineBuffer_565;
    end
    if (sel) begin
      lineBuffer_567 <= lineBuffer_566;
    end
    if (sel) begin
      lineBuffer_568 <= lineBuffer_567;
    end
    if (sel) begin
      lineBuffer_569 <= lineBuffer_568;
    end
    if (sel) begin
      lineBuffer_570 <= lineBuffer_569;
    end
    if (sel) begin
      lineBuffer_571 <= lineBuffer_570;
    end
    if (sel) begin
      lineBuffer_572 <= lineBuffer_571;
    end
    if (sel) begin
      lineBuffer_573 <= lineBuffer_572;
    end
    if (sel) begin
      lineBuffer_574 <= lineBuffer_573;
    end
    if (sel) begin
      lineBuffer_575 <= lineBuffer_574;
    end
    if (sel) begin
      lineBuffer_576 <= lineBuffer_575;
    end
    if (sel) begin
      lineBuffer_577 <= lineBuffer_576;
    end
    if (sel) begin
      lineBuffer_578 <= lineBuffer_577;
    end
    if (sel) begin
      lineBuffer_579 <= lineBuffer_578;
    end
    if (sel) begin
      lineBuffer_580 <= lineBuffer_579;
    end
    if (sel) begin
      lineBuffer_581 <= lineBuffer_580;
    end
    if (sel) begin
      lineBuffer_582 <= lineBuffer_581;
    end
    if (sel) begin
      lineBuffer_583 <= lineBuffer_582;
    end
    if (sel) begin
      lineBuffer_584 <= lineBuffer_583;
    end
    if (sel) begin
      lineBuffer_585 <= lineBuffer_584;
    end
    if (sel) begin
      lineBuffer_586 <= lineBuffer_585;
    end
    if (sel) begin
      lineBuffer_587 <= lineBuffer_586;
    end
    if (sel) begin
      lineBuffer_588 <= lineBuffer_587;
    end
    if (sel) begin
      lineBuffer_589 <= lineBuffer_588;
    end
    if (sel) begin
      lineBuffer_590 <= lineBuffer_589;
    end
    if (sel) begin
      lineBuffer_591 <= lineBuffer_590;
    end
    if (sel) begin
      lineBuffer_592 <= lineBuffer_591;
    end
    if (sel) begin
      lineBuffer_593 <= lineBuffer_592;
    end
    if (sel) begin
      lineBuffer_594 <= lineBuffer_593;
    end
    if (sel) begin
      lineBuffer_595 <= lineBuffer_594;
    end
    if (sel) begin
      lineBuffer_596 <= lineBuffer_595;
    end
    if (sel) begin
      lineBuffer_597 <= lineBuffer_596;
    end
    if (sel) begin
      lineBuffer_598 <= lineBuffer_597;
    end
    if (sel) begin
      lineBuffer_599 <= lineBuffer_598;
    end
    if (sel) begin
      lineBuffer_600 <= lineBuffer_599;
    end
    if (sel) begin
      lineBuffer_601 <= lineBuffer_600;
    end
    if (sel) begin
      lineBuffer_602 <= lineBuffer_601;
    end
    if (sel) begin
      lineBuffer_603 <= lineBuffer_602;
    end
    if (sel) begin
      lineBuffer_604 <= lineBuffer_603;
    end
    if (sel) begin
      lineBuffer_605 <= lineBuffer_604;
    end
    if (sel) begin
      lineBuffer_606 <= lineBuffer_605;
    end
    if (sel) begin
      lineBuffer_607 <= lineBuffer_606;
    end
    if (sel) begin
      lineBuffer_608 <= lineBuffer_607;
    end
    if (sel) begin
      lineBuffer_609 <= lineBuffer_608;
    end
    if (sel) begin
      lineBuffer_610 <= lineBuffer_609;
    end
    if (sel) begin
      lineBuffer_611 <= lineBuffer_610;
    end
    if (sel) begin
      lineBuffer_612 <= lineBuffer_611;
    end
    if (sel) begin
      lineBuffer_613 <= lineBuffer_612;
    end
    if (sel) begin
      lineBuffer_614 <= lineBuffer_613;
    end
    if (sel) begin
      lineBuffer_615 <= lineBuffer_614;
    end
    if (sel) begin
      lineBuffer_616 <= lineBuffer_615;
    end
    if (sel) begin
      lineBuffer_617 <= lineBuffer_616;
    end
    if (sel) begin
      lineBuffer_618 <= lineBuffer_617;
    end
    if (sel) begin
      lineBuffer_619 <= lineBuffer_618;
    end
    if (sel) begin
      lineBuffer_620 <= lineBuffer_619;
    end
    if (sel) begin
      lineBuffer_621 <= lineBuffer_620;
    end
    if (sel) begin
      lineBuffer_622 <= lineBuffer_621;
    end
    if (sel) begin
      lineBuffer_623 <= lineBuffer_622;
    end
    if (sel) begin
      lineBuffer_624 <= lineBuffer_623;
    end
    if (sel) begin
      lineBuffer_625 <= lineBuffer_624;
    end
    if (sel) begin
      lineBuffer_626 <= lineBuffer_625;
    end
    if (sel) begin
      lineBuffer_627 <= lineBuffer_626;
    end
    if (sel) begin
      lineBuffer_628 <= lineBuffer_627;
    end
    if (sel) begin
      lineBuffer_629 <= lineBuffer_628;
    end
    if (sel) begin
      lineBuffer_630 <= lineBuffer_629;
    end
    if (sel) begin
      lineBuffer_631 <= lineBuffer_630;
    end
    if (sel) begin
      lineBuffer_632 <= lineBuffer_631;
    end
    if (sel) begin
      lineBuffer_633 <= lineBuffer_632;
    end
    if (sel) begin
      lineBuffer_634 <= lineBuffer_633;
    end
    if (sel) begin
      lineBuffer_635 <= lineBuffer_634;
    end
    if (sel) begin
      lineBuffer_636 <= lineBuffer_635;
    end
    if (sel) begin
      lineBuffer_637 <= lineBuffer_636;
    end
    if (sel) begin
      lineBuffer_638 <= lineBuffer_637;
    end
    if (sel) begin
      lineBuffer_639 <= lineBuffer_638;
    end
    if (sel) begin
      lineBuffer_640 <= lineBuffer_639;
    end
    if (sel) begin
      lineBuffer_641 <= lineBuffer_640;
    end
    if (sel) begin
      lineBuffer_642 <= lineBuffer_641;
    end
    if (sel) begin
      lineBuffer_643 <= lineBuffer_642;
    end
    if (sel) begin
      lineBuffer_644 <= lineBuffer_643;
    end
    if (sel) begin
      lineBuffer_645 <= lineBuffer_644;
    end
    if (sel) begin
      lineBuffer_646 <= lineBuffer_645;
    end
    if (sel) begin
      lineBuffer_647 <= lineBuffer_646;
    end
    if (sel) begin
      lineBuffer_648 <= lineBuffer_647;
    end
    if (sel) begin
      lineBuffer_649 <= lineBuffer_648;
    end
    if (sel) begin
      lineBuffer_650 <= lineBuffer_649;
    end
    if (sel) begin
      lineBuffer_651 <= lineBuffer_650;
    end
    if (sel) begin
      lineBuffer_652 <= lineBuffer_651;
    end
    if (sel) begin
      lineBuffer_653 <= lineBuffer_652;
    end
    if (sel) begin
      lineBuffer_654 <= lineBuffer_653;
    end
    if (sel) begin
      lineBuffer_655 <= lineBuffer_654;
    end
    if (sel) begin
      lineBuffer_656 <= lineBuffer_655;
    end
    if (sel) begin
      lineBuffer_657 <= lineBuffer_656;
    end
    if (sel) begin
      lineBuffer_658 <= lineBuffer_657;
    end
    if (sel) begin
      lineBuffer_659 <= lineBuffer_658;
    end
    if (sel) begin
      lineBuffer_660 <= lineBuffer_659;
    end
    if (sel) begin
      lineBuffer_661 <= lineBuffer_660;
    end
    if (sel) begin
      lineBuffer_662 <= lineBuffer_661;
    end
    if (sel) begin
      lineBuffer_663 <= lineBuffer_662;
    end
    if (sel) begin
      lineBuffer_664 <= lineBuffer_663;
    end
    if (sel) begin
      lineBuffer_665 <= lineBuffer_664;
    end
    if (sel) begin
      lineBuffer_666 <= lineBuffer_665;
    end
    if (sel) begin
      lineBuffer_667 <= lineBuffer_666;
    end
    if (sel) begin
      lineBuffer_668 <= lineBuffer_667;
    end
    if (sel) begin
      lineBuffer_669 <= lineBuffer_668;
    end
    if (sel) begin
      lineBuffer_670 <= lineBuffer_669;
    end
    if (sel) begin
      lineBuffer_671 <= lineBuffer_670;
    end
    if (sel) begin
      lineBuffer_672 <= lineBuffer_671;
    end
    if (sel) begin
      lineBuffer_673 <= lineBuffer_672;
    end
    if (sel) begin
      lineBuffer_674 <= lineBuffer_673;
    end
    if (sel) begin
      lineBuffer_675 <= lineBuffer_674;
    end
    if (sel) begin
      lineBuffer_676 <= lineBuffer_675;
    end
    if (sel) begin
      lineBuffer_677 <= lineBuffer_676;
    end
    if (sel) begin
      lineBuffer_678 <= lineBuffer_677;
    end
    if (sel) begin
      lineBuffer_679 <= lineBuffer_678;
    end
    if (sel) begin
      lineBuffer_680 <= lineBuffer_679;
    end
    if (sel) begin
      lineBuffer_681 <= lineBuffer_680;
    end
    if (sel) begin
      lineBuffer_682 <= lineBuffer_681;
    end
    if (sel) begin
      lineBuffer_683 <= lineBuffer_682;
    end
    if (sel) begin
      lineBuffer_684 <= lineBuffer_683;
    end
    if (sel) begin
      lineBuffer_685 <= lineBuffer_684;
    end
    if (sel) begin
      lineBuffer_686 <= lineBuffer_685;
    end
    if (sel) begin
      lineBuffer_687 <= lineBuffer_686;
    end
    if (sel) begin
      lineBuffer_688 <= lineBuffer_687;
    end
    if (sel) begin
      lineBuffer_689 <= lineBuffer_688;
    end
    if (sel) begin
      lineBuffer_690 <= lineBuffer_689;
    end
    if (sel) begin
      lineBuffer_691 <= lineBuffer_690;
    end
    if (sel) begin
      lineBuffer_692 <= lineBuffer_691;
    end
    if (sel) begin
      lineBuffer_693 <= lineBuffer_692;
    end
    if (sel) begin
      lineBuffer_694 <= lineBuffer_693;
    end
    if (sel) begin
      lineBuffer_695 <= lineBuffer_694;
    end
    if (sel) begin
      lineBuffer_696 <= lineBuffer_695;
    end
    if (sel) begin
      lineBuffer_697 <= lineBuffer_696;
    end
    if (sel) begin
      lineBuffer_698 <= lineBuffer_697;
    end
    if (sel) begin
      lineBuffer_699 <= lineBuffer_698;
    end
    if (sel) begin
      lineBuffer_700 <= lineBuffer_699;
    end
    if (sel) begin
      lineBuffer_701 <= lineBuffer_700;
    end
    if (sel) begin
      lineBuffer_702 <= lineBuffer_701;
    end
    if (sel) begin
      lineBuffer_703 <= lineBuffer_702;
    end
    if (sel) begin
      lineBuffer_704 <= lineBuffer_703;
    end
    if (sel) begin
      lineBuffer_705 <= lineBuffer_704;
    end
    if (sel) begin
      lineBuffer_706 <= lineBuffer_705;
    end
    if (sel) begin
      lineBuffer_707 <= lineBuffer_706;
    end
    if (sel) begin
      lineBuffer_708 <= lineBuffer_707;
    end
    if (sel) begin
      lineBuffer_709 <= lineBuffer_708;
    end
    if (sel) begin
      lineBuffer_710 <= lineBuffer_709;
    end
    if (sel) begin
      lineBuffer_711 <= lineBuffer_710;
    end
    if (sel) begin
      lineBuffer_712 <= lineBuffer_711;
    end
    if (sel) begin
      lineBuffer_713 <= lineBuffer_712;
    end
    if (sel) begin
      lineBuffer_714 <= lineBuffer_713;
    end
    if (sel) begin
      lineBuffer_715 <= lineBuffer_714;
    end
    if (sel) begin
      lineBuffer_716 <= lineBuffer_715;
    end
    if (sel) begin
      lineBuffer_717 <= lineBuffer_716;
    end
    if (sel) begin
      lineBuffer_718 <= lineBuffer_717;
    end
    if (sel) begin
      lineBuffer_719 <= lineBuffer_718;
    end
    if (sel) begin
      lineBuffer_720 <= lineBuffer_719;
    end
    if (sel) begin
      lineBuffer_721 <= lineBuffer_720;
    end
    if (sel) begin
      lineBuffer_722 <= lineBuffer_721;
    end
    if (sel) begin
      lineBuffer_723 <= lineBuffer_722;
    end
    if (sel) begin
      lineBuffer_724 <= lineBuffer_723;
    end
    if (sel) begin
      lineBuffer_725 <= lineBuffer_724;
    end
    if (sel) begin
      lineBuffer_726 <= lineBuffer_725;
    end
    if (sel) begin
      lineBuffer_727 <= lineBuffer_726;
    end
    if (sel) begin
      lineBuffer_728 <= lineBuffer_727;
    end
    if (sel) begin
      lineBuffer_729 <= lineBuffer_728;
    end
    if (sel) begin
      lineBuffer_730 <= lineBuffer_729;
    end
    if (sel) begin
      lineBuffer_731 <= lineBuffer_730;
    end
    if (sel) begin
      lineBuffer_732 <= lineBuffer_731;
    end
    if (sel) begin
      lineBuffer_733 <= lineBuffer_732;
    end
    if (sel) begin
      lineBuffer_734 <= lineBuffer_733;
    end
    if (sel) begin
      lineBuffer_735 <= lineBuffer_734;
    end
    if (sel) begin
      lineBuffer_736 <= lineBuffer_735;
    end
    if (sel) begin
      lineBuffer_737 <= lineBuffer_736;
    end
    if (sel) begin
      lineBuffer_738 <= lineBuffer_737;
    end
    if (sel) begin
      lineBuffer_739 <= lineBuffer_738;
    end
    if (sel) begin
      lineBuffer_740 <= lineBuffer_739;
    end
    if (sel) begin
      lineBuffer_741 <= lineBuffer_740;
    end
    if (sel) begin
      lineBuffer_742 <= lineBuffer_741;
    end
    if (sel) begin
      lineBuffer_743 <= lineBuffer_742;
    end
    if (sel) begin
      lineBuffer_744 <= lineBuffer_743;
    end
    if (sel) begin
      lineBuffer_745 <= lineBuffer_744;
    end
    if (sel) begin
      lineBuffer_746 <= lineBuffer_745;
    end
    if (sel) begin
      lineBuffer_747 <= lineBuffer_746;
    end
    if (sel) begin
      lineBuffer_748 <= lineBuffer_747;
    end
    if (sel) begin
      lineBuffer_749 <= lineBuffer_748;
    end
    if (sel) begin
      lineBuffer_750 <= lineBuffer_749;
    end
    if (sel) begin
      lineBuffer_751 <= lineBuffer_750;
    end
    if (sel) begin
      lineBuffer_752 <= lineBuffer_751;
    end
    if (sel) begin
      lineBuffer_753 <= lineBuffer_752;
    end
    if (sel) begin
      lineBuffer_754 <= lineBuffer_753;
    end
    if (sel) begin
      lineBuffer_755 <= lineBuffer_754;
    end
    if (sel) begin
      lineBuffer_756 <= lineBuffer_755;
    end
    if (sel) begin
      lineBuffer_757 <= lineBuffer_756;
    end
    if (sel) begin
      lineBuffer_758 <= lineBuffer_757;
    end
    if (sel) begin
      lineBuffer_759 <= lineBuffer_758;
    end
    if (sel) begin
      lineBuffer_760 <= lineBuffer_759;
    end
    if (sel) begin
      lineBuffer_761 <= lineBuffer_760;
    end
    if (sel) begin
      lineBuffer_762 <= lineBuffer_761;
    end
    if (sel) begin
      lineBuffer_763 <= lineBuffer_762;
    end
    if (sel) begin
      lineBuffer_764 <= lineBuffer_763;
    end
    if (sel) begin
      lineBuffer_765 <= lineBuffer_764;
    end
    if (sel) begin
      lineBuffer_766 <= lineBuffer_765;
    end
    if (sel) begin
      lineBuffer_767 <= lineBuffer_766;
    end
    if (sel) begin
      windowBuffer_0 <= windowBuffer_1;
    end
    if (sel) begin
      windowBuffer_1 <= windowBuffer_2;
    end
    if (sel) begin
      windowBuffer_2 <= _T_797;
    end
    if (sel) begin
      windowBuffer_3 <= windowBuffer_4;
    end
    if (sel) begin
      windowBuffer_4 <= windowBuffer_5;
    end
    if (sel) begin
      windowBuffer_5 <= _T_801;
    end
    if (sel) begin
      windowBuffer_6 <= windowBuffer_7;
    end
    if (sel) begin
      windowBuffer_7 <= windowBuffer_8;
    end
    if (sel) begin
      windowBuffer_8 <= _T_805;
    end
  end
endmodule
module NonMaxSupression(
  input        clock,
  input        reset,
  output       io_enq_ready,
  input        io_enq_valid,
  input  [1:0] io_enq_bits_grad_dir,
  input  [7:0] io_enq_bits_value,
  input        io_enq_user,
  input        io_enq_last,
  input        io_deq_ready,
  output       io_deq_valid,
  output [7:0] io_deq_bits,
  output       io_deq_user,
  output       io_deq_last
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
  reg [31:0] _RAND_64;
  reg [31:0] _RAND_65;
  reg [31:0] _RAND_66;
  reg [31:0] _RAND_67;
  reg [31:0] _RAND_68;
  reg [31:0] _RAND_69;
  reg [31:0] _RAND_70;
  reg [31:0] _RAND_71;
  reg [31:0] _RAND_72;
  reg [31:0] _RAND_73;
  reg [31:0] _RAND_74;
  reg [31:0] _RAND_75;
  reg [31:0] _RAND_76;
  reg [31:0] _RAND_77;
  reg [31:0] _RAND_78;
  reg [31:0] _RAND_79;
  reg [31:0] _RAND_80;
  reg [31:0] _RAND_81;
  reg [31:0] _RAND_82;
  reg [31:0] _RAND_83;
  reg [31:0] _RAND_84;
  reg [31:0] _RAND_85;
  reg [31:0] _RAND_86;
  reg [31:0] _RAND_87;
  reg [31:0] _RAND_88;
  reg [31:0] _RAND_89;
  reg [31:0] _RAND_90;
  reg [31:0] _RAND_91;
  reg [31:0] _RAND_92;
  reg [31:0] _RAND_93;
  reg [31:0] _RAND_94;
  reg [31:0] _RAND_95;
  reg [31:0] _RAND_96;
  reg [31:0] _RAND_97;
  reg [31:0] _RAND_98;
  reg [31:0] _RAND_99;
  reg [31:0] _RAND_100;
  reg [31:0] _RAND_101;
  reg [31:0] _RAND_102;
  reg [31:0] _RAND_103;
  reg [31:0] _RAND_104;
  reg [31:0] _RAND_105;
  reg [31:0] _RAND_106;
  reg [31:0] _RAND_107;
  reg [31:0] _RAND_108;
  reg [31:0] _RAND_109;
  reg [31:0] _RAND_110;
  reg [31:0] _RAND_111;
  reg [31:0] _RAND_112;
  reg [31:0] _RAND_113;
  reg [31:0] _RAND_114;
  reg [31:0] _RAND_115;
  reg [31:0] _RAND_116;
  reg [31:0] _RAND_117;
  reg [31:0] _RAND_118;
  reg [31:0] _RAND_119;
  reg [31:0] _RAND_120;
  reg [31:0] _RAND_121;
  reg [31:0] _RAND_122;
  reg [31:0] _RAND_123;
  reg [31:0] _RAND_124;
  reg [31:0] _RAND_125;
  reg [31:0] _RAND_126;
  reg [31:0] _RAND_127;
  reg [31:0] _RAND_128;
  reg [31:0] _RAND_129;
  reg [31:0] _RAND_130;
  reg [31:0] _RAND_131;
  reg [31:0] _RAND_132;
  reg [31:0] _RAND_133;
  reg [31:0] _RAND_134;
  reg [31:0] _RAND_135;
  reg [31:0] _RAND_136;
  reg [31:0] _RAND_137;
  reg [31:0] _RAND_138;
  reg [31:0] _RAND_139;
  reg [31:0] _RAND_140;
  reg [31:0] _RAND_141;
  reg [31:0] _RAND_142;
  reg [31:0] _RAND_143;
  reg [31:0] _RAND_144;
  reg [31:0] _RAND_145;
  reg [31:0] _RAND_146;
  reg [31:0] _RAND_147;
  reg [31:0] _RAND_148;
  reg [31:0] _RAND_149;
  reg [31:0] _RAND_150;
  reg [31:0] _RAND_151;
  reg [31:0] _RAND_152;
  reg [31:0] _RAND_153;
  reg [31:0] _RAND_154;
  reg [31:0] _RAND_155;
  reg [31:0] _RAND_156;
  reg [31:0] _RAND_157;
  reg [31:0] _RAND_158;
  reg [31:0] _RAND_159;
  reg [31:0] _RAND_160;
  reg [31:0] _RAND_161;
  reg [31:0] _RAND_162;
  reg [31:0] _RAND_163;
  reg [31:0] _RAND_164;
  reg [31:0] _RAND_165;
  reg [31:0] _RAND_166;
  reg [31:0] _RAND_167;
  reg [31:0] _RAND_168;
  reg [31:0] _RAND_169;
  reg [31:0] _RAND_170;
  reg [31:0] _RAND_171;
  reg [31:0] _RAND_172;
  reg [31:0] _RAND_173;
  reg [31:0] _RAND_174;
  reg [31:0] _RAND_175;
  reg [31:0] _RAND_176;
  reg [31:0] _RAND_177;
  reg [31:0] _RAND_178;
  reg [31:0] _RAND_179;
  reg [31:0] _RAND_180;
  reg [31:0] _RAND_181;
  reg [31:0] _RAND_182;
  reg [31:0] _RAND_183;
  reg [31:0] _RAND_184;
  reg [31:0] _RAND_185;
  reg [31:0] _RAND_186;
  reg [31:0] _RAND_187;
  reg [31:0] _RAND_188;
  reg [31:0] _RAND_189;
  reg [31:0] _RAND_190;
  reg [31:0] _RAND_191;
  reg [31:0] _RAND_192;
  reg [31:0] _RAND_193;
  reg [31:0] _RAND_194;
  reg [31:0] _RAND_195;
  reg [31:0] _RAND_196;
  reg [31:0] _RAND_197;
  reg [31:0] _RAND_198;
  reg [31:0] _RAND_199;
  reg [31:0] _RAND_200;
  reg [31:0] _RAND_201;
  reg [31:0] _RAND_202;
  reg [31:0] _RAND_203;
  reg [31:0] _RAND_204;
  reg [31:0] _RAND_205;
  reg [31:0] _RAND_206;
  reg [31:0] _RAND_207;
  reg [31:0] _RAND_208;
  reg [31:0] _RAND_209;
  reg [31:0] _RAND_210;
  reg [31:0] _RAND_211;
  reg [31:0] _RAND_212;
  reg [31:0] _RAND_213;
  reg [31:0] _RAND_214;
  reg [31:0] _RAND_215;
  reg [31:0] _RAND_216;
  reg [31:0] _RAND_217;
  reg [31:0] _RAND_218;
  reg [31:0] _RAND_219;
  reg [31:0] _RAND_220;
  reg [31:0] _RAND_221;
  reg [31:0] _RAND_222;
  reg [31:0] _RAND_223;
  reg [31:0] _RAND_224;
  reg [31:0] _RAND_225;
  reg [31:0] _RAND_226;
  reg [31:0] _RAND_227;
  reg [31:0] _RAND_228;
  reg [31:0] _RAND_229;
  reg [31:0] _RAND_230;
  reg [31:0] _RAND_231;
  reg [31:0] _RAND_232;
  reg [31:0] _RAND_233;
  reg [31:0] _RAND_234;
  reg [31:0] _RAND_235;
  reg [31:0] _RAND_236;
  reg [31:0] _RAND_237;
  reg [31:0] _RAND_238;
  reg [31:0] _RAND_239;
  reg [31:0] _RAND_240;
  reg [31:0] _RAND_241;
  reg [31:0] _RAND_242;
  reg [31:0] _RAND_243;
  reg [31:0] _RAND_244;
  reg [31:0] _RAND_245;
  reg [31:0] _RAND_246;
  reg [31:0] _RAND_247;
  reg [31:0] _RAND_248;
  reg [31:0] _RAND_249;
  reg [31:0] _RAND_250;
  reg [31:0] _RAND_251;
  reg [31:0] _RAND_252;
  reg [31:0] _RAND_253;
  reg [31:0] _RAND_254;
  reg [31:0] _RAND_255;
  reg [31:0] _RAND_256;
  reg [31:0] _RAND_257;
  reg [31:0] _RAND_258;
  reg [31:0] _RAND_259;
  reg [31:0] _RAND_260;
  reg [31:0] _RAND_261;
  reg [31:0] _RAND_262;
  reg [31:0] _RAND_263;
  reg [31:0] _RAND_264;
  reg [31:0] _RAND_265;
  reg [31:0] _RAND_266;
  reg [31:0] _RAND_267;
  reg [31:0] _RAND_268;
  reg [31:0] _RAND_269;
  reg [31:0] _RAND_270;
  reg [31:0] _RAND_271;
  reg [31:0] _RAND_272;
  reg [31:0] _RAND_273;
  reg [31:0] _RAND_274;
  reg [31:0] _RAND_275;
  reg [31:0] _RAND_276;
  reg [31:0] _RAND_277;
  reg [31:0] _RAND_278;
  reg [31:0] _RAND_279;
  reg [31:0] _RAND_280;
  reg [31:0] _RAND_281;
  reg [31:0] _RAND_282;
  reg [31:0] _RAND_283;
  reg [31:0] _RAND_284;
  reg [31:0] _RAND_285;
  reg [31:0] _RAND_286;
  reg [31:0] _RAND_287;
  reg [31:0] _RAND_288;
  reg [31:0] _RAND_289;
  reg [31:0] _RAND_290;
  reg [31:0] _RAND_291;
  reg [31:0] _RAND_292;
  reg [31:0] _RAND_293;
  reg [31:0] _RAND_294;
  reg [31:0] _RAND_295;
  reg [31:0] _RAND_296;
  reg [31:0] _RAND_297;
  reg [31:0] _RAND_298;
  reg [31:0] _RAND_299;
  reg [31:0] _RAND_300;
  reg [31:0] _RAND_301;
  reg [31:0] _RAND_302;
  reg [31:0] _RAND_303;
  reg [31:0] _RAND_304;
  reg [31:0] _RAND_305;
  reg [31:0] _RAND_306;
  reg [31:0] _RAND_307;
  reg [31:0] _RAND_308;
  reg [31:0] _RAND_309;
  reg [31:0] _RAND_310;
  reg [31:0] _RAND_311;
  reg [31:0] _RAND_312;
  reg [31:0] _RAND_313;
  reg [31:0] _RAND_314;
  reg [31:0] _RAND_315;
  reg [31:0] _RAND_316;
  reg [31:0] _RAND_317;
  reg [31:0] _RAND_318;
  reg [31:0] _RAND_319;
  reg [31:0] _RAND_320;
  reg [31:0] _RAND_321;
  reg [31:0] _RAND_322;
  reg [31:0] _RAND_323;
  reg [31:0] _RAND_324;
  reg [31:0] _RAND_325;
  reg [31:0] _RAND_326;
  reg [31:0] _RAND_327;
  reg [31:0] _RAND_328;
  reg [31:0] _RAND_329;
  reg [31:0] _RAND_330;
  reg [31:0] _RAND_331;
  reg [31:0] _RAND_332;
  reg [31:0] _RAND_333;
  reg [31:0] _RAND_334;
  reg [31:0] _RAND_335;
  reg [31:0] _RAND_336;
  reg [31:0] _RAND_337;
  reg [31:0] _RAND_338;
  reg [31:0] _RAND_339;
  reg [31:0] _RAND_340;
  reg [31:0] _RAND_341;
  reg [31:0] _RAND_342;
  reg [31:0] _RAND_343;
  reg [31:0] _RAND_344;
  reg [31:0] _RAND_345;
  reg [31:0] _RAND_346;
  reg [31:0] _RAND_347;
  reg [31:0] _RAND_348;
  reg [31:0] _RAND_349;
  reg [31:0] _RAND_350;
  reg [31:0] _RAND_351;
  reg [31:0] _RAND_352;
  reg [31:0] _RAND_353;
  reg [31:0] _RAND_354;
  reg [31:0] _RAND_355;
  reg [31:0] _RAND_356;
  reg [31:0] _RAND_357;
  reg [31:0] _RAND_358;
  reg [31:0] _RAND_359;
  reg [31:0] _RAND_360;
  reg [31:0] _RAND_361;
  reg [31:0] _RAND_362;
  reg [31:0] _RAND_363;
  reg [31:0] _RAND_364;
  reg [31:0] _RAND_365;
  reg [31:0] _RAND_366;
  reg [31:0] _RAND_367;
  reg [31:0] _RAND_368;
  reg [31:0] _RAND_369;
  reg [31:0] _RAND_370;
  reg [31:0] _RAND_371;
  reg [31:0] _RAND_372;
  reg [31:0] _RAND_373;
  reg [31:0] _RAND_374;
  reg [31:0] _RAND_375;
  reg [31:0] _RAND_376;
  reg [31:0] _RAND_377;
  reg [31:0] _RAND_378;
  reg [31:0] _RAND_379;
  reg [31:0] _RAND_380;
  reg [31:0] _RAND_381;
  reg [31:0] _RAND_382;
  reg [31:0] _RAND_383;
  reg [31:0] _RAND_384;
  reg [31:0] _RAND_385;
  reg [31:0] _RAND_386;
  reg [31:0] _RAND_387;
  reg [31:0] _RAND_388;
  reg [31:0] _RAND_389;
  reg [31:0] _RAND_390;
  reg [31:0] _RAND_391;
  reg [31:0] _RAND_392;
  reg [31:0] _RAND_393;
  reg [31:0] _RAND_394;
  reg [31:0] _RAND_395;
  reg [31:0] _RAND_396;
  reg [31:0] _RAND_397;
  reg [31:0] _RAND_398;
  reg [31:0] _RAND_399;
  reg [31:0] _RAND_400;
  reg [31:0] _RAND_401;
  reg [31:0] _RAND_402;
  reg [31:0] _RAND_403;
  reg [31:0] _RAND_404;
  reg [31:0] _RAND_405;
  reg [31:0] _RAND_406;
  reg [31:0] _RAND_407;
  reg [31:0] _RAND_408;
  reg [31:0] _RAND_409;
  reg [31:0] _RAND_410;
  reg [31:0] _RAND_411;
  reg [31:0] _RAND_412;
  reg [31:0] _RAND_413;
  reg [31:0] _RAND_414;
  reg [31:0] _RAND_415;
  reg [31:0] _RAND_416;
  reg [31:0] _RAND_417;
  reg [31:0] _RAND_418;
  reg [31:0] _RAND_419;
  reg [31:0] _RAND_420;
  reg [31:0] _RAND_421;
  reg [31:0] _RAND_422;
  reg [31:0] _RAND_423;
  reg [31:0] _RAND_424;
  reg [31:0] _RAND_425;
  reg [31:0] _RAND_426;
  reg [31:0] _RAND_427;
  reg [31:0] _RAND_428;
  reg [31:0] _RAND_429;
  reg [31:0] _RAND_430;
  reg [31:0] _RAND_431;
  reg [31:0] _RAND_432;
  reg [31:0] _RAND_433;
  reg [31:0] _RAND_434;
  reg [31:0] _RAND_435;
  reg [31:0] _RAND_436;
  reg [31:0] _RAND_437;
  reg [31:0] _RAND_438;
  reg [31:0] _RAND_439;
  reg [31:0] _RAND_440;
  reg [31:0] _RAND_441;
  reg [31:0] _RAND_442;
  reg [31:0] _RAND_443;
  reg [31:0] _RAND_444;
  reg [31:0] _RAND_445;
  reg [31:0] _RAND_446;
  reg [31:0] _RAND_447;
  reg [31:0] _RAND_448;
  reg [31:0] _RAND_449;
  reg [31:0] _RAND_450;
  reg [31:0] _RAND_451;
  reg [31:0] _RAND_452;
  reg [31:0] _RAND_453;
  reg [31:0] _RAND_454;
  reg [31:0] _RAND_455;
  reg [31:0] _RAND_456;
  reg [31:0] _RAND_457;
  reg [31:0] _RAND_458;
  reg [31:0] _RAND_459;
  reg [31:0] _RAND_460;
  reg [31:0] _RAND_461;
  reg [31:0] _RAND_462;
  reg [31:0] _RAND_463;
  reg [31:0] _RAND_464;
  reg [31:0] _RAND_465;
  reg [31:0] _RAND_466;
  reg [31:0] _RAND_467;
  reg [31:0] _RAND_468;
  reg [31:0] _RAND_469;
  reg [31:0] _RAND_470;
  reg [31:0] _RAND_471;
  reg [31:0] _RAND_472;
  reg [31:0] _RAND_473;
  reg [31:0] _RAND_474;
  reg [31:0] _RAND_475;
  reg [31:0] _RAND_476;
  reg [31:0] _RAND_477;
  reg [31:0] _RAND_478;
  reg [31:0] _RAND_479;
  reg [31:0] _RAND_480;
  reg [31:0] _RAND_481;
  reg [31:0] _RAND_482;
  reg [31:0] _RAND_483;
  reg [31:0] _RAND_484;
  reg [31:0] _RAND_485;
  reg [31:0] _RAND_486;
  reg [31:0] _RAND_487;
  reg [31:0] _RAND_488;
  reg [31:0] _RAND_489;
  reg [31:0] _RAND_490;
  reg [31:0] _RAND_491;
  reg [31:0] _RAND_492;
  reg [31:0] _RAND_493;
  reg [31:0] _RAND_494;
  reg [31:0] _RAND_495;
  reg [31:0] _RAND_496;
  reg [31:0] _RAND_497;
  reg [31:0] _RAND_498;
  reg [31:0] _RAND_499;
  reg [31:0] _RAND_500;
  reg [31:0] _RAND_501;
  reg [31:0] _RAND_502;
  reg [31:0] _RAND_503;
  reg [31:0] _RAND_504;
  reg [31:0] _RAND_505;
  reg [31:0] _RAND_506;
  reg [31:0] _RAND_507;
  reg [31:0] _RAND_508;
  reg [31:0] _RAND_509;
  reg [31:0] _RAND_510;
  reg [31:0] _RAND_511;
  reg [31:0] _RAND_512;
  reg [31:0] _RAND_513;
  reg [31:0] _RAND_514;
  reg [31:0] _RAND_515;
  reg [31:0] _RAND_516;
  reg [31:0] _RAND_517;
  reg [31:0] _RAND_518;
  reg [31:0] _RAND_519;
  reg [31:0] _RAND_520;
  reg [31:0] _RAND_521;
  reg [31:0] _RAND_522;
  reg [31:0] _RAND_523;
  reg [31:0] _RAND_524;
  reg [31:0] _RAND_525;
  reg [31:0] _RAND_526;
  reg [31:0] _RAND_527;
  reg [31:0] _RAND_528;
  reg [31:0] _RAND_529;
  reg [31:0] _RAND_530;
  reg [31:0] _RAND_531;
  reg [31:0] _RAND_532;
  reg [31:0] _RAND_533;
  reg [31:0] _RAND_534;
  reg [31:0] _RAND_535;
  reg [31:0] _RAND_536;
  reg [31:0] _RAND_537;
  reg [31:0] _RAND_538;
  reg [31:0] _RAND_539;
  reg [31:0] _RAND_540;
  reg [31:0] _RAND_541;
  reg [31:0] _RAND_542;
  reg [31:0] _RAND_543;
  reg [31:0] _RAND_544;
  reg [31:0] _RAND_545;
  reg [31:0] _RAND_546;
  reg [31:0] _RAND_547;
  reg [31:0] _RAND_548;
  reg [31:0] _RAND_549;
  reg [31:0] _RAND_550;
  reg [31:0] _RAND_551;
  reg [31:0] _RAND_552;
  reg [31:0] _RAND_553;
  reg [31:0] _RAND_554;
  reg [31:0] _RAND_555;
  reg [31:0] _RAND_556;
  reg [31:0] _RAND_557;
  reg [31:0] _RAND_558;
  reg [31:0] _RAND_559;
  reg [31:0] _RAND_560;
  reg [31:0] _RAND_561;
  reg [31:0] _RAND_562;
  reg [31:0] _RAND_563;
  reg [31:0] _RAND_564;
  reg [31:0] _RAND_565;
  reg [31:0] _RAND_566;
  reg [31:0] _RAND_567;
  reg [31:0] _RAND_568;
  reg [31:0] _RAND_569;
  reg [31:0] _RAND_570;
  reg [31:0] _RAND_571;
  reg [31:0] _RAND_572;
  reg [31:0] _RAND_573;
  reg [31:0] _RAND_574;
  reg [31:0] _RAND_575;
  reg [31:0] _RAND_576;
  reg [31:0] _RAND_577;
  reg [31:0] _RAND_578;
  reg [31:0] _RAND_579;
  reg [31:0] _RAND_580;
  reg [31:0] _RAND_581;
  reg [31:0] _RAND_582;
  reg [31:0] _RAND_583;
  reg [31:0] _RAND_584;
  reg [31:0] _RAND_585;
  reg [31:0] _RAND_586;
  reg [31:0] _RAND_587;
  reg [31:0] _RAND_588;
  reg [31:0] _RAND_589;
  reg [31:0] _RAND_590;
  reg [31:0] _RAND_591;
  reg [31:0] _RAND_592;
  reg [31:0] _RAND_593;
  reg [31:0] _RAND_594;
  reg [31:0] _RAND_595;
  reg [31:0] _RAND_596;
  reg [31:0] _RAND_597;
  reg [31:0] _RAND_598;
  reg [31:0] _RAND_599;
  reg [31:0] _RAND_600;
  reg [31:0] _RAND_601;
  reg [31:0] _RAND_602;
  reg [31:0] _RAND_603;
  reg [31:0] _RAND_604;
  reg [31:0] _RAND_605;
  reg [31:0] _RAND_606;
  reg [31:0] _RAND_607;
  reg [31:0] _RAND_608;
  reg [31:0] _RAND_609;
  reg [31:0] _RAND_610;
  reg [31:0] _RAND_611;
  reg [31:0] _RAND_612;
  reg [31:0] _RAND_613;
  reg [31:0] _RAND_614;
  reg [31:0] _RAND_615;
  reg [31:0] _RAND_616;
  reg [31:0] _RAND_617;
  reg [31:0] _RAND_618;
  reg [31:0] _RAND_619;
  reg [31:0] _RAND_620;
  reg [31:0] _RAND_621;
  reg [31:0] _RAND_622;
  reg [31:0] _RAND_623;
  reg [31:0] _RAND_624;
  reg [31:0] _RAND_625;
  reg [31:0] _RAND_626;
  reg [31:0] _RAND_627;
  reg [31:0] _RAND_628;
  reg [31:0] _RAND_629;
  reg [31:0] _RAND_630;
  reg [31:0] _RAND_631;
  reg [31:0] _RAND_632;
  reg [31:0] _RAND_633;
  reg [31:0] _RAND_634;
  reg [31:0] _RAND_635;
  reg [31:0] _RAND_636;
  reg [31:0] _RAND_637;
  reg [31:0] _RAND_638;
  reg [31:0] _RAND_639;
  reg [31:0] _RAND_640;
  reg [31:0] _RAND_641;
  reg [31:0] _RAND_642;
  reg [31:0] _RAND_643;
  reg [31:0] _RAND_644;
  reg [31:0] _RAND_645;
  reg [31:0] _RAND_646;
  reg [31:0] _RAND_647;
  reg [31:0] _RAND_648;
  reg [31:0] _RAND_649;
  reg [31:0] _RAND_650;
  reg [31:0] _RAND_651;
  reg [31:0] _RAND_652;
  reg [31:0] _RAND_653;
  reg [31:0] _RAND_654;
  reg [31:0] _RAND_655;
  reg [31:0] _RAND_656;
  reg [31:0] _RAND_657;
  reg [31:0] _RAND_658;
  reg [31:0] _RAND_659;
  reg [31:0] _RAND_660;
  reg [31:0] _RAND_661;
  reg [31:0] _RAND_662;
  reg [31:0] _RAND_663;
  reg [31:0] _RAND_664;
  reg [31:0] _RAND_665;
  reg [31:0] _RAND_666;
  reg [31:0] _RAND_667;
  reg [31:0] _RAND_668;
  reg [31:0] _RAND_669;
  reg [31:0] _RAND_670;
  reg [31:0] _RAND_671;
  reg [31:0] _RAND_672;
  reg [31:0] _RAND_673;
  reg [31:0] _RAND_674;
  reg [31:0] _RAND_675;
  reg [31:0] _RAND_676;
  reg [31:0] _RAND_677;
  reg [31:0] _RAND_678;
  reg [31:0] _RAND_679;
  reg [31:0] _RAND_680;
  reg [31:0] _RAND_681;
  reg [31:0] _RAND_682;
  reg [31:0] _RAND_683;
  reg [31:0] _RAND_684;
  reg [31:0] _RAND_685;
  reg [31:0] _RAND_686;
  reg [31:0] _RAND_687;
  reg [31:0] _RAND_688;
  reg [31:0] _RAND_689;
  reg [31:0] _RAND_690;
  reg [31:0] _RAND_691;
  reg [31:0] _RAND_692;
  reg [31:0] _RAND_693;
  reg [31:0] _RAND_694;
  reg [31:0] _RAND_695;
  reg [31:0] _RAND_696;
  reg [31:0] _RAND_697;
  reg [31:0] _RAND_698;
  reg [31:0] _RAND_699;
  reg [31:0] _RAND_700;
  reg [31:0] _RAND_701;
  reg [31:0] _RAND_702;
  reg [31:0] _RAND_703;
  reg [31:0] _RAND_704;
  reg [31:0] _RAND_705;
  reg [31:0] _RAND_706;
  reg [31:0] _RAND_707;
  reg [31:0] _RAND_708;
  reg [31:0] _RAND_709;
  reg [31:0] _RAND_710;
  reg [31:0] _RAND_711;
  reg [31:0] _RAND_712;
  reg [31:0] _RAND_713;
  reg [31:0] _RAND_714;
  reg [31:0] _RAND_715;
  reg [31:0] _RAND_716;
  reg [31:0] _RAND_717;
  reg [31:0] _RAND_718;
  reg [31:0] _RAND_719;
  reg [31:0] _RAND_720;
  reg [31:0] _RAND_721;
  reg [31:0] _RAND_722;
  reg [31:0] _RAND_723;
  reg [31:0] _RAND_724;
  reg [31:0] _RAND_725;
  reg [31:0] _RAND_726;
  reg [31:0] _RAND_727;
  reg [31:0] _RAND_728;
  reg [31:0] _RAND_729;
  reg [31:0] _RAND_730;
  reg [31:0] _RAND_731;
  reg [31:0] _RAND_732;
  reg [31:0] _RAND_733;
  reg [31:0] _RAND_734;
  reg [31:0] _RAND_735;
  reg [31:0] _RAND_736;
  reg [31:0] _RAND_737;
  reg [31:0] _RAND_738;
  reg [31:0] _RAND_739;
  reg [31:0] _RAND_740;
  reg [31:0] _RAND_741;
  reg [31:0] _RAND_742;
  reg [31:0] _RAND_743;
  reg [31:0] _RAND_744;
  reg [31:0] _RAND_745;
  reg [31:0] _RAND_746;
  reg [31:0] _RAND_747;
  reg [31:0] _RAND_748;
  reg [31:0] _RAND_749;
  reg [31:0] _RAND_750;
  reg [31:0] _RAND_751;
  reg [31:0] _RAND_752;
  reg [31:0] _RAND_753;
  reg [31:0] _RAND_754;
  reg [31:0] _RAND_755;
  reg [31:0] _RAND_756;
  reg [31:0] _RAND_757;
  reg [31:0] _RAND_758;
  reg [31:0] _RAND_759;
  reg [31:0] _RAND_760;
  reg [31:0] _RAND_761;
  reg [31:0] _RAND_762;
  reg [31:0] _RAND_763;
  reg [31:0] _RAND_764;
  reg [31:0] _RAND_765;
  reg [31:0] _RAND_766;
  reg [31:0] _RAND_767;
  reg [31:0] _RAND_768;
  reg [31:0] _RAND_769;
  reg [31:0] _RAND_770;
  reg [31:0] _RAND_771;
  reg [31:0] _RAND_772;
  reg [31:0] _RAND_773;
  reg [31:0] _RAND_774;
  reg [31:0] _RAND_775;
  reg [31:0] _RAND_776;
  reg [31:0] _RAND_777;
  reg [31:0] _RAND_778;
  reg [31:0] _RAND_779;
  reg [31:0] _RAND_780;
  reg [31:0] _RAND_781;
  reg [31:0] _RAND_782;
  reg [31:0] _RAND_783;
  reg [31:0] _RAND_784;
  reg [31:0] _RAND_785;
  reg [31:0] _RAND_786;
  reg [31:0] _RAND_787;
  reg [31:0] _RAND_788;
  reg [31:0] _RAND_789;
  reg [31:0] _RAND_790;
  reg [31:0] _RAND_791;
  reg [31:0] _RAND_792;
  reg [31:0] _RAND_793;
  reg [31:0] _RAND_794;
  reg [31:0] _RAND_795;
  reg [31:0] _RAND_796;
  reg [31:0] _RAND_797;
  reg [31:0] _RAND_798;
  reg [31:0] _RAND_799;
  reg [31:0] _RAND_800;
  reg [31:0] _RAND_801;
  reg [31:0] _RAND_802;
  reg [31:0] _RAND_803;
  reg [31:0] _RAND_804;
  reg [31:0] _RAND_805;
  reg [31:0] _RAND_806;
  reg [31:0] _RAND_807;
  reg [31:0] _RAND_808;
  reg [31:0] _RAND_809;
  reg [31:0] _RAND_810;
  reg [31:0] _RAND_811;
  reg [31:0] _RAND_812;
  reg [31:0] _RAND_813;
  reg [31:0] _RAND_814;
  reg [31:0] _RAND_815;
  reg [31:0] _RAND_816;
  reg [31:0] _RAND_817;
  reg [31:0] _RAND_818;
  reg [31:0] _RAND_819;
  reg [31:0] _RAND_820;
  reg [31:0] _RAND_821;
  reg [31:0] _RAND_822;
  reg [31:0] _RAND_823;
  reg [31:0] _RAND_824;
  reg [31:0] _RAND_825;
  reg [31:0] _RAND_826;
  reg [31:0] _RAND_827;
  reg [31:0] _RAND_828;
  reg [31:0] _RAND_829;
  reg [31:0] _RAND_830;
  reg [31:0] _RAND_831;
  reg [31:0] _RAND_832;
  reg [31:0] _RAND_833;
  reg [31:0] _RAND_834;
  reg [31:0] _RAND_835;
  reg [31:0] _RAND_836;
  reg [31:0] _RAND_837;
  reg [31:0] _RAND_838;
  reg [31:0] _RAND_839;
  reg [31:0] _RAND_840;
  reg [31:0] _RAND_841;
  reg [31:0] _RAND_842;
  reg [31:0] _RAND_843;
  reg [31:0] _RAND_844;
  reg [31:0] _RAND_845;
  reg [31:0] _RAND_846;
  reg [31:0] _RAND_847;
  reg [31:0] _RAND_848;
  reg [31:0] _RAND_849;
  reg [31:0] _RAND_850;
  reg [31:0] _RAND_851;
  reg [31:0] _RAND_852;
  reg [31:0] _RAND_853;
  reg [31:0] _RAND_854;
  reg [31:0] _RAND_855;
  reg [31:0] _RAND_856;
  reg [31:0] _RAND_857;
  reg [31:0] _RAND_858;
  reg [31:0] _RAND_859;
  reg [31:0] _RAND_860;
  reg [31:0] _RAND_861;
  reg [31:0] _RAND_862;
  reg [31:0] _RAND_863;
  reg [31:0] _RAND_864;
  reg [31:0] _RAND_865;
  reg [31:0] _RAND_866;
  reg [31:0] _RAND_867;
  reg [31:0] _RAND_868;
  reg [31:0] _RAND_869;
  reg [31:0] _RAND_870;
  reg [31:0] _RAND_871;
  reg [31:0] _RAND_872;
  reg [31:0] _RAND_873;
  reg [31:0] _RAND_874;
  reg [31:0] _RAND_875;
  reg [31:0] _RAND_876;
  reg [31:0] _RAND_877;
  reg [31:0] _RAND_878;
  reg [31:0] _RAND_879;
  reg [31:0] _RAND_880;
  reg [31:0] _RAND_881;
  reg [31:0] _RAND_882;
  reg [31:0] _RAND_883;
  reg [31:0] _RAND_884;
  reg [31:0] _RAND_885;
  reg [31:0] _RAND_886;
  reg [31:0] _RAND_887;
  reg [31:0] _RAND_888;
  reg [31:0] _RAND_889;
  reg [31:0] _RAND_890;
  reg [31:0] _RAND_891;
  reg [31:0] _RAND_892;
  reg [31:0] _RAND_893;
  reg [31:0] _RAND_894;
  reg [31:0] _RAND_895;
  reg [31:0] _RAND_896;
  reg [31:0] _RAND_897;
  reg [31:0] _RAND_898;
  reg [31:0] _RAND_899;
  reg [31:0] _RAND_900;
  reg [31:0] _RAND_901;
  reg [31:0] _RAND_902;
  reg [31:0] _RAND_903;
  reg [31:0] _RAND_904;
  reg [31:0] _RAND_905;
  reg [31:0] _RAND_906;
  reg [31:0] _RAND_907;
  reg [31:0] _RAND_908;
  reg [31:0] _RAND_909;
  reg [31:0] _RAND_910;
  reg [31:0] _RAND_911;
  reg [31:0] _RAND_912;
  reg [31:0] _RAND_913;
  reg [31:0] _RAND_914;
  reg [31:0] _RAND_915;
  reg [31:0] _RAND_916;
  reg [31:0] _RAND_917;
  reg [31:0] _RAND_918;
  reg [31:0] _RAND_919;
  reg [31:0] _RAND_920;
  reg [31:0] _RAND_921;
  reg [31:0] _RAND_922;
  reg [31:0] _RAND_923;
  reg [31:0] _RAND_924;
  reg [31:0] _RAND_925;
  reg [31:0] _RAND_926;
  reg [31:0] _RAND_927;
  reg [31:0] _RAND_928;
  reg [31:0] _RAND_929;
  reg [31:0] _RAND_930;
  reg [31:0] _RAND_931;
  reg [31:0] _RAND_932;
  reg [31:0] _RAND_933;
  reg [31:0] _RAND_934;
  reg [31:0] _RAND_935;
  reg [31:0] _RAND_936;
  reg [31:0] _RAND_937;
  reg [31:0] _RAND_938;
  reg [31:0] _RAND_939;
  reg [31:0] _RAND_940;
  reg [31:0] _RAND_941;
  reg [31:0] _RAND_942;
  reg [31:0] _RAND_943;
  reg [31:0] _RAND_944;
  reg [31:0] _RAND_945;
  reg [31:0] _RAND_946;
  reg [31:0] _RAND_947;
  reg [31:0] _RAND_948;
  reg [31:0] _RAND_949;
  reg [31:0] _RAND_950;
  reg [31:0] _RAND_951;
  reg [31:0] _RAND_952;
  reg [31:0] _RAND_953;
  reg [31:0] _RAND_954;
  reg [31:0] _RAND_955;
  reg [31:0] _RAND_956;
  reg [31:0] _RAND_957;
  reg [31:0] _RAND_958;
  reg [31:0] _RAND_959;
  reg [31:0] _RAND_960;
  reg [31:0] _RAND_961;
  reg [31:0] _RAND_962;
  reg [31:0] _RAND_963;
  reg [31:0] _RAND_964;
  reg [31:0] _RAND_965;
  reg [31:0] _RAND_966;
  reg [31:0] _RAND_967;
  reg [31:0] _RAND_968;
  reg [31:0] _RAND_969;
  reg [31:0] _RAND_970;
  reg [31:0] _RAND_971;
  reg [31:0] _RAND_972;
  reg [31:0] _RAND_973;
  reg [31:0] _RAND_974;
  reg [31:0] _RAND_975;
  reg [31:0] _RAND_976;
  reg [31:0] _RAND_977;
  reg [31:0] _RAND_978;
  reg [31:0] _RAND_979;
  reg [31:0] _RAND_980;
  reg [31:0] _RAND_981;
  reg [31:0] _RAND_982;
  reg [31:0] _RAND_983;
  reg [31:0] _RAND_984;
  reg [31:0] _RAND_985;
  reg [31:0] _RAND_986;
  reg [31:0] _RAND_987;
  reg [31:0] _RAND_988;
  reg [31:0] _RAND_989;
  reg [31:0] _RAND_990;
  reg [31:0] _RAND_991;
  reg [31:0] _RAND_992;
  reg [31:0] _RAND_993;
  reg [31:0] _RAND_994;
  reg [31:0] _RAND_995;
  reg [31:0] _RAND_996;
  reg [31:0] _RAND_997;
  reg [31:0] _RAND_998;
  reg [31:0] _RAND_999;
  reg [31:0] _RAND_1000;
  reg [31:0] _RAND_1001;
  reg [31:0] _RAND_1002;
  reg [31:0] _RAND_1003;
  reg [31:0] _RAND_1004;
  reg [31:0] _RAND_1005;
  reg [31:0] _RAND_1006;
  reg [31:0] _RAND_1007;
  reg [31:0] _RAND_1008;
  reg [31:0] _RAND_1009;
  reg [31:0] _RAND_1010;
  reg [31:0] _RAND_1011;
  reg [31:0] _RAND_1012;
  reg [31:0] _RAND_1013;
  reg [31:0] _RAND_1014;
  reg [31:0] _RAND_1015;
  reg [31:0] _RAND_1016;
  reg [31:0] _RAND_1017;
  reg [31:0] _RAND_1018;
  reg [31:0] _RAND_1019;
  reg [31:0] _RAND_1020;
  reg [31:0] _RAND_1021;
  reg [31:0] _RAND_1022;
  reg [31:0] _RAND_1023;
  reg [31:0] _RAND_1024;
  reg [31:0] _RAND_1025;
  reg [31:0] _RAND_1026;
  reg [31:0] _RAND_1027;
  reg [31:0] _RAND_1028;
  reg [31:0] _RAND_1029;
  reg [31:0] _RAND_1030;
  reg [31:0] _RAND_1031;
  reg [31:0] _RAND_1032;
  reg [31:0] _RAND_1033;
  reg [31:0] _RAND_1034;
  reg [31:0] _RAND_1035;
  reg [31:0] _RAND_1036;
  reg [31:0] _RAND_1037;
  reg [31:0] _RAND_1038;
  reg [31:0] _RAND_1039;
  reg [31:0] _RAND_1040;
  reg [31:0] _RAND_1041;
  reg [31:0] _RAND_1042;
  reg [31:0] _RAND_1043;
  reg [31:0] _RAND_1044;
  reg [31:0] _RAND_1045;
  reg [31:0] _RAND_1046;
  reg [31:0] _RAND_1047;
  reg [31:0] _RAND_1048;
  reg [31:0] _RAND_1049;
  reg [31:0] _RAND_1050;
  reg [31:0] _RAND_1051;
  reg [31:0] _RAND_1052;
  reg [31:0] _RAND_1053;
  reg [31:0] _RAND_1054;
  reg [31:0] _RAND_1055;
  reg [31:0] _RAND_1056;
  reg [31:0] _RAND_1057;
  reg [31:0] _RAND_1058;
  reg [31:0] _RAND_1059;
  reg [31:0] _RAND_1060;
  reg [31:0] _RAND_1061;
  reg [31:0] _RAND_1062;
  reg [31:0] _RAND_1063;
  reg [31:0] _RAND_1064;
  reg [31:0] _RAND_1065;
  reg [31:0] _RAND_1066;
  reg [31:0] _RAND_1067;
  reg [31:0] _RAND_1068;
  reg [31:0] _RAND_1069;
  reg [31:0] _RAND_1070;
  reg [31:0] _RAND_1071;
  reg [31:0] _RAND_1072;
  reg [31:0] _RAND_1073;
  reg [31:0] _RAND_1074;
  reg [31:0] _RAND_1075;
  reg [31:0] _RAND_1076;
  reg [31:0] _RAND_1077;
  reg [31:0] _RAND_1078;
  reg [31:0] _RAND_1079;
  reg [31:0] _RAND_1080;
  reg [31:0] _RAND_1081;
  reg [31:0] _RAND_1082;
  reg [31:0] _RAND_1083;
  reg [31:0] _RAND_1084;
  reg [31:0] _RAND_1085;
  reg [31:0] _RAND_1086;
  reg [31:0] _RAND_1087;
  reg [31:0] _RAND_1088;
  reg [31:0] _RAND_1089;
  reg [31:0] _RAND_1090;
  reg [31:0] _RAND_1091;
  reg [31:0] _RAND_1092;
  reg [31:0] _RAND_1093;
  reg [31:0] _RAND_1094;
  reg [31:0] _RAND_1095;
  reg [31:0] _RAND_1096;
  reg [31:0] _RAND_1097;
  reg [31:0] _RAND_1098;
  reg [31:0] _RAND_1099;
  reg [31:0] _RAND_1100;
  reg [31:0] _RAND_1101;
  reg [31:0] _RAND_1102;
  reg [31:0] _RAND_1103;
  reg [31:0] _RAND_1104;
  reg [31:0] _RAND_1105;
  reg [31:0] _RAND_1106;
  reg [31:0] _RAND_1107;
  reg [31:0] _RAND_1108;
  reg [31:0] _RAND_1109;
  reg [31:0] _RAND_1110;
  reg [31:0] _RAND_1111;
  reg [31:0] _RAND_1112;
  reg [31:0] _RAND_1113;
  reg [31:0] _RAND_1114;
  reg [31:0] _RAND_1115;
  reg [31:0] _RAND_1116;
  reg [31:0] _RAND_1117;
  reg [31:0] _RAND_1118;
  reg [31:0] _RAND_1119;
  reg [31:0] _RAND_1120;
  reg [31:0] _RAND_1121;
  reg [31:0] _RAND_1122;
  reg [31:0] _RAND_1123;
  reg [31:0] _RAND_1124;
  reg [31:0] _RAND_1125;
  reg [31:0] _RAND_1126;
  reg [31:0] _RAND_1127;
  reg [31:0] _RAND_1128;
  reg [31:0] _RAND_1129;
  reg [31:0] _RAND_1130;
  reg [31:0] _RAND_1131;
  reg [31:0] _RAND_1132;
  reg [31:0] _RAND_1133;
  reg [31:0] _RAND_1134;
  reg [31:0] _RAND_1135;
  reg [31:0] _RAND_1136;
  reg [31:0] _RAND_1137;
  reg [31:0] _RAND_1138;
  reg [31:0] _RAND_1139;
  reg [31:0] _RAND_1140;
  reg [31:0] _RAND_1141;
  reg [31:0] _RAND_1142;
  reg [31:0] _RAND_1143;
  reg [31:0] _RAND_1144;
  reg [31:0] _RAND_1145;
  reg [31:0] _RAND_1146;
  reg [31:0] _RAND_1147;
  reg [31:0] _RAND_1148;
  reg [31:0] _RAND_1149;
  reg [31:0] _RAND_1150;
  reg [31:0] _RAND_1151;
  reg [31:0] _RAND_1152;
  reg [31:0] _RAND_1153;
  reg [31:0] _RAND_1154;
  reg [31:0] _RAND_1155;
  reg [31:0] _RAND_1156;
  reg [31:0] _RAND_1157;
  reg [31:0] _RAND_1158;
  reg [31:0] _RAND_1159;
  reg [31:0] _RAND_1160;
  reg [31:0] _RAND_1161;
  reg [31:0] _RAND_1162;
  reg [31:0] _RAND_1163;
  reg [31:0] _RAND_1164;
  reg [31:0] _RAND_1165;
  reg [31:0] _RAND_1166;
  reg [31:0] _RAND_1167;
  reg [31:0] _RAND_1168;
  reg [31:0] _RAND_1169;
  reg [31:0] _RAND_1170;
  reg [31:0] _RAND_1171;
  reg [31:0] _RAND_1172;
  reg [31:0] _RAND_1173;
  reg [31:0] _RAND_1174;
  reg [31:0] _RAND_1175;
  reg [31:0] _RAND_1176;
  reg [31:0] _RAND_1177;
  reg [31:0] _RAND_1178;
  reg [31:0] _RAND_1179;
  reg [31:0] _RAND_1180;
  reg [31:0] _RAND_1181;
  reg [31:0] _RAND_1182;
  reg [31:0] _RAND_1183;
  reg [31:0] _RAND_1184;
  reg [31:0] _RAND_1185;
  reg [31:0] _RAND_1186;
  reg [31:0] _RAND_1187;
  reg [31:0] _RAND_1188;
  reg [31:0] _RAND_1189;
  reg [31:0] _RAND_1190;
  reg [31:0] _RAND_1191;
  reg [31:0] _RAND_1192;
  reg [31:0] _RAND_1193;
  reg [31:0] _RAND_1194;
  reg [31:0] _RAND_1195;
  reg [31:0] _RAND_1196;
  reg [31:0] _RAND_1197;
  reg [31:0] _RAND_1198;
  reg [31:0] _RAND_1199;
  reg [31:0] _RAND_1200;
  reg [31:0] _RAND_1201;
  reg [31:0] _RAND_1202;
  reg [31:0] _RAND_1203;
  reg [31:0] _RAND_1204;
  reg [31:0] _RAND_1205;
  reg [31:0] _RAND_1206;
  reg [31:0] _RAND_1207;
  reg [31:0] _RAND_1208;
  reg [31:0] _RAND_1209;
  reg [31:0] _RAND_1210;
  reg [31:0] _RAND_1211;
  reg [31:0] _RAND_1212;
  reg [31:0] _RAND_1213;
  reg [31:0] _RAND_1214;
  reg [31:0] _RAND_1215;
  reg [31:0] _RAND_1216;
  reg [31:0] _RAND_1217;
  reg [31:0] _RAND_1218;
  reg [31:0] _RAND_1219;
  reg [31:0] _RAND_1220;
  reg [31:0] _RAND_1221;
  reg [31:0] _RAND_1222;
  reg [31:0] _RAND_1223;
  reg [31:0] _RAND_1224;
  reg [31:0] _RAND_1225;
  reg [31:0] _RAND_1226;
  reg [31:0] _RAND_1227;
  reg [31:0] _RAND_1228;
  reg [31:0] _RAND_1229;
  reg [31:0] _RAND_1230;
  reg [31:0] _RAND_1231;
  reg [31:0] _RAND_1232;
  reg [31:0] _RAND_1233;
  reg [31:0] _RAND_1234;
  reg [31:0] _RAND_1235;
  reg [31:0] _RAND_1236;
  reg [31:0] _RAND_1237;
  reg [31:0] _RAND_1238;
  reg [31:0] _RAND_1239;
  reg [31:0] _RAND_1240;
  reg [31:0] _RAND_1241;
  reg [31:0] _RAND_1242;
  reg [31:0] _RAND_1243;
  reg [31:0] _RAND_1244;
  reg [31:0] _RAND_1245;
  reg [31:0] _RAND_1246;
  reg [31:0] _RAND_1247;
  reg [31:0] _RAND_1248;
  reg [31:0] _RAND_1249;
  reg [31:0] _RAND_1250;
  reg [31:0] _RAND_1251;
  reg [31:0] _RAND_1252;
  reg [31:0] _RAND_1253;
  reg [31:0] _RAND_1254;
  reg [31:0] _RAND_1255;
  reg [31:0] _RAND_1256;
  reg [31:0] _RAND_1257;
  reg [31:0] _RAND_1258;
  reg [31:0] _RAND_1259;
  reg [31:0] _RAND_1260;
  reg [31:0] _RAND_1261;
  reg [31:0] _RAND_1262;
  reg [31:0] _RAND_1263;
  reg [31:0] _RAND_1264;
  reg [31:0] _RAND_1265;
  reg [31:0] _RAND_1266;
  reg [31:0] _RAND_1267;
  reg [31:0] _RAND_1268;
  reg [31:0] _RAND_1269;
  reg [31:0] _RAND_1270;
  reg [31:0] _RAND_1271;
  reg [31:0] _RAND_1272;
  reg [31:0] _RAND_1273;
  reg [31:0] _RAND_1274;
  reg [31:0] _RAND_1275;
  reg [31:0] _RAND_1276;
  reg [31:0] _RAND_1277;
  reg [31:0] _RAND_1278;
  reg [31:0] _RAND_1279;
  reg [31:0] _RAND_1280;
  reg [31:0] _RAND_1281;
  reg [31:0] _RAND_1282;
  reg [31:0] _RAND_1283;
  reg [31:0] _RAND_1284;
  reg [31:0] _RAND_1285;
  reg [31:0] _RAND_1286;
  reg [31:0] _RAND_1287;
  reg [31:0] _RAND_1288;
  reg [31:0] _RAND_1289;
  reg [31:0] _RAND_1290;
  reg [31:0] _RAND_1291;
  reg [31:0] _RAND_1292;
  reg [31:0] _RAND_1293;
  reg [31:0] _RAND_1294;
  reg [31:0] _RAND_1295;
  reg [31:0] _RAND_1296;
  reg [31:0] _RAND_1297;
  reg [31:0] _RAND_1298;
  reg [31:0] _RAND_1299;
`endif // RANDOMIZE_REG_INIT
  reg [1:0] stateReg; // @[ChiselImProc.scala 62:28]
  reg [1:0] dataReg_grad_dir; // @[ChiselImProc.scala 64:23]
  reg [7:0] dataReg_value; // @[ChiselImProc.scala 64:23]
  reg [1:0] shadowReg_grad_dir; // @[ChiselImProc.scala 66:25]
  reg [7:0] shadowReg_value; // @[ChiselImProc.scala 66:25]
  reg  userReg; // @[ChiselImProc.scala 67:23]
  reg  shadowUserReg; // @[ChiselImProc.scala 68:29]
  reg  lastReg; // @[ChiselImProc.scala 69:23]
  reg  shadowLastReg; // @[ChiselImProc.scala 70:29]
  reg [1:0] lineBuffer_0_grad_dir; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_0_value; // @[ChiselImProc.scala 346:25]
  reg [1:0] lineBuffer_1_grad_dir; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_1_value; // @[ChiselImProc.scala 346:25]
  reg [1:0] lineBuffer_2_grad_dir; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_2_value; // @[ChiselImProc.scala 346:25]
  reg [1:0] lineBuffer_3_grad_dir; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_3_value; // @[ChiselImProc.scala 346:25]
  reg [1:0] lineBuffer_4_grad_dir; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_4_value; // @[ChiselImProc.scala 346:25]
  reg [1:0] lineBuffer_5_grad_dir; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_5_value; // @[ChiselImProc.scala 346:25]
  reg [1:0] lineBuffer_6_grad_dir; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_6_value; // @[ChiselImProc.scala 346:25]
  reg [1:0] lineBuffer_7_grad_dir; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_7_value; // @[ChiselImProc.scala 346:25]
  reg [1:0] lineBuffer_8_grad_dir; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_8_value; // @[ChiselImProc.scala 346:25]
  reg [1:0] lineBuffer_9_grad_dir; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_9_value; // @[ChiselImProc.scala 346:25]
  reg [1:0] lineBuffer_10_grad_dir; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_10_value; // @[ChiselImProc.scala 346:25]
  reg [1:0] lineBuffer_11_grad_dir; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_11_value; // @[ChiselImProc.scala 346:25]
  reg [1:0] lineBuffer_12_grad_dir; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_12_value; // @[ChiselImProc.scala 346:25]
  reg [1:0] lineBuffer_13_grad_dir; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_13_value; // @[ChiselImProc.scala 346:25]
  reg [1:0] lineBuffer_14_grad_dir; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_14_value; // @[ChiselImProc.scala 346:25]
  reg [1:0] lineBuffer_15_grad_dir; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_15_value; // @[ChiselImProc.scala 346:25]
  reg [1:0] lineBuffer_16_grad_dir; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_16_value; // @[ChiselImProc.scala 346:25]
  reg [1:0] lineBuffer_17_grad_dir; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_17_value; // @[ChiselImProc.scala 346:25]
  reg [1:0] lineBuffer_18_grad_dir; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_18_value; // @[ChiselImProc.scala 346:25]
  reg [1:0] lineBuffer_19_grad_dir; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_19_value; // @[ChiselImProc.scala 346:25]
  reg [1:0] lineBuffer_20_grad_dir; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_20_value; // @[ChiselImProc.scala 346:25]
  reg [1:0] lineBuffer_21_grad_dir; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_21_value; // @[ChiselImProc.scala 346:25]
  reg [1:0] lineBuffer_22_grad_dir; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_22_value; // @[ChiselImProc.scala 346:25]
  reg [1:0] lineBuffer_23_grad_dir; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_23_value; // @[ChiselImProc.scala 346:25]
  reg [1:0] lineBuffer_24_grad_dir; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_24_value; // @[ChiselImProc.scala 346:25]
  reg [1:0] lineBuffer_25_grad_dir; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_25_value; // @[ChiselImProc.scala 346:25]
  reg [1:0] lineBuffer_26_grad_dir; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_26_value; // @[ChiselImProc.scala 346:25]
  reg [1:0] lineBuffer_27_grad_dir; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_27_value; // @[ChiselImProc.scala 346:25]
  reg [1:0] lineBuffer_28_grad_dir; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_28_value; // @[ChiselImProc.scala 346:25]
  reg [1:0] lineBuffer_29_grad_dir; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_29_value; // @[ChiselImProc.scala 346:25]
  reg [1:0] lineBuffer_30_grad_dir; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_30_value; // @[ChiselImProc.scala 346:25]
  reg [1:0] lineBuffer_31_grad_dir; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_31_value; // @[ChiselImProc.scala 346:25]
  reg [1:0] lineBuffer_32_grad_dir; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_32_value; // @[ChiselImProc.scala 346:25]
  reg [1:0] lineBuffer_33_grad_dir; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_33_value; // @[ChiselImProc.scala 346:25]
  reg [1:0] lineBuffer_34_grad_dir; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_34_value; // @[ChiselImProc.scala 346:25]
  reg [1:0] lineBuffer_35_grad_dir; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_35_value; // @[ChiselImProc.scala 346:25]
  reg [1:0] lineBuffer_36_grad_dir; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_36_value; // @[ChiselImProc.scala 346:25]
  reg [1:0] lineBuffer_37_grad_dir; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_37_value; // @[ChiselImProc.scala 346:25]
  reg [1:0] lineBuffer_38_grad_dir; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_38_value; // @[ChiselImProc.scala 346:25]
  reg [1:0] lineBuffer_39_grad_dir; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_39_value; // @[ChiselImProc.scala 346:25]
  reg [1:0] lineBuffer_40_grad_dir; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_40_value; // @[ChiselImProc.scala 346:25]
  reg [1:0] lineBuffer_41_grad_dir; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_41_value; // @[ChiselImProc.scala 346:25]
  reg [1:0] lineBuffer_42_grad_dir; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_42_value; // @[ChiselImProc.scala 346:25]
  reg [1:0] lineBuffer_43_grad_dir; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_43_value; // @[ChiselImProc.scala 346:25]
  reg [1:0] lineBuffer_44_grad_dir; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_44_value; // @[ChiselImProc.scala 346:25]
  reg [1:0] lineBuffer_45_grad_dir; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_45_value; // @[ChiselImProc.scala 346:25]
  reg [1:0] lineBuffer_46_grad_dir; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_46_value; // @[ChiselImProc.scala 346:25]
  reg [1:0] lineBuffer_47_grad_dir; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_47_value; // @[ChiselImProc.scala 346:25]
  reg [1:0] lineBuffer_48_grad_dir; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_48_value; // @[ChiselImProc.scala 346:25]
  reg [1:0] lineBuffer_49_grad_dir; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_49_value; // @[ChiselImProc.scala 346:25]
  reg [1:0] lineBuffer_50_grad_dir; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_50_value; // @[ChiselImProc.scala 346:25]
  reg [1:0] lineBuffer_51_grad_dir; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_51_value; // @[ChiselImProc.scala 346:25]
  reg [1:0] lineBuffer_52_grad_dir; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_52_value; // @[ChiselImProc.scala 346:25]
  reg [1:0] lineBuffer_53_grad_dir; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_53_value; // @[ChiselImProc.scala 346:25]
  reg [1:0] lineBuffer_54_grad_dir; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_54_value; // @[ChiselImProc.scala 346:25]
  reg [1:0] lineBuffer_55_grad_dir; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_55_value; // @[ChiselImProc.scala 346:25]
  reg [1:0] lineBuffer_56_grad_dir; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_56_value; // @[ChiselImProc.scala 346:25]
  reg [1:0] lineBuffer_57_grad_dir; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_57_value; // @[ChiselImProc.scala 346:25]
  reg [1:0] lineBuffer_58_grad_dir; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_58_value; // @[ChiselImProc.scala 346:25]
  reg [1:0] lineBuffer_59_grad_dir; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_59_value; // @[ChiselImProc.scala 346:25]
  reg [1:0] lineBuffer_60_grad_dir; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_60_value; // @[ChiselImProc.scala 346:25]
  reg [1:0] lineBuffer_61_grad_dir; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_61_value; // @[ChiselImProc.scala 346:25]
  reg [1:0] lineBuffer_62_grad_dir; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_62_value; // @[ChiselImProc.scala 346:25]
  reg [1:0] lineBuffer_63_grad_dir; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_63_value; // @[ChiselImProc.scala 346:25]
  reg [1:0] lineBuffer_64_grad_dir; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_64_value; // @[ChiselImProc.scala 346:25]
  reg [1:0] lineBuffer_65_grad_dir; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_65_value; // @[ChiselImProc.scala 346:25]
  reg [1:0] lineBuffer_66_grad_dir; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_66_value; // @[ChiselImProc.scala 346:25]
  reg [1:0] lineBuffer_67_grad_dir; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_67_value; // @[ChiselImProc.scala 346:25]
  reg [1:0] lineBuffer_68_grad_dir; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_68_value; // @[ChiselImProc.scala 346:25]
  reg [1:0] lineBuffer_69_grad_dir; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_69_value; // @[ChiselImProc.scala 346:25]
  reg [1:0] lineBuffer_70_grad_dir; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_70_value; // @[ChiselImProc.scala 346:25]
  reg [1:0] lineBuffer_71_grad_dir; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_71_value; // @[ChiselImProc.scala 346:25]
  reg [1:0] lineBuffer_72_grad_dir; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_72_value; // @[ChiselImProc.scala 346:25]
  reg [1:0] lineBuffer_73_grad_dir; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_73_value; // @[ChiselImProc.scala 346:25]
  reg [1:0] lineBuffer_74_grad_dir; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_74_value; // @[ChiselImProc.scala 346:25]
  reg [1:0] lineBuffer_75_grad_dir; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_75_value; // @[ChiselImProc.scala 346:25]
  reg [1:0] lineBuffer_76_grad_dir; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_76_value; // @[ChiselImProc.scala 346:25]
  reg [1:0] lineBuffer_77_grad_dir; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_77_value; // @[ChiselImProc.scala 346:25]
  reg [1:0] lineBuffer_78_grad_dir; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_78_value; // @[ChiselImProc.scala 346:25]
  reg [1:0] lineBuffer_79_grad_dir; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_79_value; // @[ChiselImProc.scala 346:25]
  reg [1:0] lineBuffer_80_grad_dir; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_80_value; // @[ChiselImProc.scala 346:25]
  reg [1:0] lineBuffer_81_grad_dir; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_81_value; // @[ChiselImProc.scala 346:25]
  reg [1:0] lineBuffer_82_grad_dir; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_82_value; // @[ChiselImProc.scala 346:25]
  reg [1:0] lineBuffer_83_grad_dir; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_83_value; // @[ChiselImProc.scala 346:25]
  reg [1:0] lineBuffer_84_grad_dir; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_84_value; // @[ChiselImProc.scala 346:25]
  reg [1:0] lineBuffer_85_grad_dir; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_85_value; // @[ChiselImProc.scala 346:25]
  reg [1:0] lineBuffer_86_grad_dir; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_86_value; // @[ChiselImProc.scala 346:25]
  reg [1:0] lineBuffer_87_grad_dir; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_87_value; // @[ChiselImProc.scala 346:25]
  reg [1:0] lineBuffer_88_grad_dir; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_88_value; // @[ChiselImProc.scala 346:25]
  reg [1:0] lineBuffer_89_grad_dir; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_89_value; // @[ChiselImProc.scala 346:25]
  reg [1:0] lineBuffer_90_grad_dir; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_90_value; // @[ChiselImProc.scala 346:25]
  reg [1:0] lineBuffer_91_grad_dir; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_91_value; // @[ChiselImProc.scala 346:25]
  reg [1:0] lineBuffer_92_grad_dir; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_92_value; // @[ChiselImProc.scala 346:25]
  reg [1:0] lineBuffer_93_grad_dir; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_93_value; // @[ChiselImProc.scala 346:25]
  reg [1:0] lineBuffer_94_grad_dir; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_94_value; // @[ChiselImProc.scala 346:25]
  reg [1:0] lineBuffer_95_grad_dir; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_95_value; // @[ChiselImProc.scala 346:25]
  reg [1:0] lineBuffer_96_grad_dir; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_96_value; // @[ChiselImProc.scala 346:25]
  reg [1:0] lineBuffer_97_grad_dir; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_97_value; // @[ChiselImProc.scala 346:25]
  reg [1:0] lineBuffer_98_grad_dir; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_98_value; // @[ChiselImProc.scala 346:25]
  reg [1:0] lineBuffer_99_grad_dir; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_99_value; // @[ChiselImProc.scala 346:25]
  reg [1:0] lineBuffer_100_grad_dir; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_100_value; // @[ChiselImProc.scala 346:25]
  reg [1:0] lineBuffer_101_grad_dir; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_101_value; // @[ChiselImProc.scala 346:25]
  reg [1:0] lineBuffer_102_grad_dir; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_102_value; // @[ChiselImProc.scala 346:25]
  reg [1:0] lineBuffer_103_grad_dir; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_103_value; // @[ChiselImProc.scala 346:25]
  reg [1:0] lineBuffer_104_grad_dir; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_104_value; // @[ChiselImProc.scala 346:25]
  reg [1:0] lineBuffer_105_grad_dir; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_105_value; // @[ChiselImProc.scala 346:25]
  reg [1:0] lineBuffer_106_grad_dir; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_106_value; // @[ChiselImProc.scala 346:25]
  reg [1:0] lineBuffer_107_grad_dir; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_107_value; // @[ChiselImProc.scala 346:25]
  reg [1:0] lineBuffer_108_grad_dir; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_108_value; // @[ChiselImProc.scala 346:25]
  reg [1:0] lineBuffer_109_grad_dir; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_109_value; // @[ChiselImProc.scala 346:25]
  reg [1:0] lineBuffer_110_grad_dir; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_110_value; // @[ChiselImProc.scala 346:25]
  reg [1:0] lineBuffer_111_grad_dir; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_111_value; // @[ChiselImProc.scala 346:25]
  reg [1:0] lineBuffer_112_grad_dir; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_112_value; // @[ChiselImProc.scala 346:25]
  reg [1:0] lineBuffer_113_grad_dir; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_113_value; // @[ChiselImProc.scala 346:25]
  reg [1:0] lineBuffer_114_grad_dir; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_114_value; // @[ChiselImProc.scala 346:25]
  reg [1:0] lineBuffer_115_grad_dir; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_115_value; // @[ChiselImProc.scala 346:25]
  reg [1:0] lineBuffer_116_grad_dir; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_116_value; // @[ChiselImProc.scala 346:25]
  reg [1:0] lineBuffer_117_grad_dir; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_117_value; // @[ChiselImProc.scala 346:25]
  reg [1:0] lineBuffer_118_grad_dir; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_118_value; // @[ChiselImProc.scala 346:25]
  reg [1:0] lineBuffer_119_grad_dir; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_119_value; // @[ChiselImProc.scala 346:25]
  reg [1:0] lineBuffer_120_grad_dir; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_120_value; // @[ChiselImProc.scala 346:25]
  reg [1:0] lineBuffer_121_grad_dir; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_121_value; // @[ChiselImProc.scala 346:25]
  reg [1:0] lineBuffer_122_grad_dir; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_122_value; // @[ChiselImProc.scala 346:25]
  reg [1:0] lineBuffer_123_grad_dir; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_123_value; // @[ChiselImProc.scala 346:25]
  reg [1:0] lineBuffer_124_grad_dir; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_124_value; // @[ChiselImProc.scala 346:25]
  reg [1:0] lineBuffer_125_grad_dir; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_125_value; // @[ChiselImProc.scala 346:25]
  reg [1:0] lineBuffer_126_grad_dir; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_126_value; // @[ChiselImProc.scala 346:25]
  reg [1:0] lineBuffer_127_grad_dir; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_127_value; // @[ChiselImProc.scala 346:25]
  reg [1:0] lineBuffer_128_grad_dir; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_128_value; // @[ChiselImProc.scala 346:25]
  reg [1:0] lineBuffer_129_grad_dir; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_129_value; // @[ChiselImProc.scala 346:25]
  reg [1:0] lineBuffer_130_grad_dir; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_130_value; // @[ChiselImProc.scala 346:25]
  reg [1:0] lineBuffer_131_grad_dir; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_131_value; // @[ChiselImProc.scala 346:25]
  reg [1:0] lineBuffer_132_grad_dir; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_132_value; // @[ChiselImProc.scala 346:25]
  reg [1:0] lineBuffer_133_grad_dir; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_133_value; // @[ChiselImProc.scala 346:25]
  reg [1:0] lineBuffer_134_grad_dir; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_134_value; // @[ChiselImProc.scala 346:25]
  reg [1:0] lineBuffer_135_grad_dir; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_135_value; // @[ChiselImProc.scala 346:25]
  reg [1:0] lineBuffer_136_grad_dir; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_136_value; // @[ChiselImProc.scala 346:25]
  reg [1:0] lineBuffer_137_grad_dir; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_137_value; // @[ChiselImProc.scala 346:25]
  reg [1:0] lineBuffer_138_grad_dir; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_138_value; // @[ChiselImProc.scala 346:25]
  reg [1:0] lineBuffer_139_grad_dir; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_139_value; // @[ChiselImProc.scala 346:25]
  reg [1:0] lineBuffer_140_grad_dir; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_140_value; // @[ChiselImProc.scala 346:25]
  reg [1:0] lineBuffer_141_grad_dir; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_141_value; // @[ChiselImProc.scala 346:25]
  reg [1:0] lineBuffer_142_grad_dir; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_142_value; // @[ChiselImProc.scala 346:25]
  reg [1:0] lineBuffer_143_grad_dir; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_143_value; // @[ChiselImProc.scala 346:25]
  reg [1:0] lineBuffer_144_grad_dir; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_144_value; // @[ChiselImProc.scala 346:25]
  reg [1:0] lineBuffer_145_grad_dir; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_145_value; // @[ChiselImProc.scala 346:25]
  reg [1:0] lineBuffer_146_grad_dir; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_146_value; // @[ChiselImProc.scala 346:25]
  reg [1:0] lineBuffer_147_grad_dir; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_147_value; // @[ChiselImProc.scala 346:25]
  reg [1:0] lineBuffer_148_grad_dir; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_148_value; // @[ChiselImProc.scala 346:25]
  reg [1:0] lineBuffer_149_grad_dir; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_149_value; // @[ChiselImProc.scala 346:25]
  reg [1:0] lineBuffer_150_grad_dir; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_150_value; // @[ChiselImProc.scala 346:25]
  reg [1:0] lineBuffer_151_grad_dir; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_151_value; // @[ChiselImProc.scala 346:25]
  reg [1:0] lineBuffer_152_grad_dir; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_152_value; // @[ChiselImProc.scala 346:25]
  reg [1:0] lineBuffer_153_grad_dir; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_153_value; // @[ChiselImProc.scala 346:25]
  reg [1:0] lineBuffer_154_grad_dir; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_154_value; // @[ChiselImProc.scala 346:25]
  reg [1:0] lineBuffer_155_grad_dir; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_155_value; // @[ChiselImProc.scala 346:25]
  reg [1:0] lineBuffer_156_grad_dir; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_156_value; // @[ChiselImProc.scala 346:25]
  reg [1:0] lineBuffer_157_grad_dir; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_157_value; // @[ChiselImProc.scala 346:25]
  reg [1:0] lineBuffer_158_grad_dir; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_158_value; // @[ChiselImProc.scala 346:25]
  reg [1:0] lineBuffer_159_grad_dir; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_159_value; // @[ChiselImProc.scala 346:25]
  reg [1:0] lineBuffer_160_grad_dir; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_160_value; // @[ChiselImProc.scala 346:25]
  reg [1:0] lineBuffer_161_grad_dir; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_161_value; // @[ChiselImProc.scala 346:25]
  reg [1:0] lineBuffer_162_grad_dir; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_162_value; // @[ChiselImProc.scala 346:25]
  reg [1:0] lineBuffer_163_grad_dir; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_163_value; // @[ChiselImProc.scala 346:25]
  reg [1:0] lineBuffer_164_grad_dir; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_164_value; // @[ChiselImProc.scala 346:25]
  reg [1:0] lineBuffer_165_grad_dir; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_165_value; // @[ChiselImProc.scala 346:25]
  reg [1:0] lineBuffer_166_grad_dir; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_166_value; // @[ChiselImProc.scala 346:25]
  reg [1:0] lineBuffer_167_grad_dir; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_167_value; // @[ChiselImProc.scala 346:25]
  reg [1:0] lineBuffer_168_grad_dir; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_168_value; // @[ChiselImProc.scala 346:25]
  reg [1:0] lineBuffer_169_grad_dir; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_169_value; // @[ChiselImProc.scala 346:25]
  reg [1:0] lineBuffer_170_grad_dir; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_170_value; // @[ChiselImProc.scala 346:25]
  reg [1:0] lineBuffer_171_grad_dir; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_171_value; // @[ChiselImProc.scala 346:25]
  reg [1:0] lineBuffer_172_grad_dir; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_172_value; // @[ChiselImProc.scala 346:25]
  reg [1:0] lineBuffer_173_grad_dir; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_173_value; // @[ChiselImProc.scala 346:25]
  reg [1:0] lineBuffer_174_grad_dir; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_174_value; // @[ChiselImProc.scala 346:25]
  reg [1:0] lineBuffer_175_grad_dir; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_175_value; // @[ChiselImProc.scala 346:25]
  reg [1:0] lineBuffer_176_grad_dir; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_176_value; // @[ChiselImProc.scala 346:25]
  reg [1:0] lineBuffer_177_grad_dir; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_177_value; // @[ChiselImProc.scala 346:25]
  reg [1:0] lineBuffer_178_grad_dir; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_178_value; // @[ChiselImProc.scala 346:25]
  reg [1:0] lineBuffer_179_grad_dir; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_179_value; // @[ChiselImProc.scala 346:25]
  reg [1:0] lineBuffer_180_grad_dir; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_180_value; // @[ChiselImProc.scala 346:25]
  reg [1:0] lineBuffer_181_grad_dir; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_181_value; // @[ChiselImProc.scala 346:25]
  reg [1:0] lineBuffer_182_grad_dir; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_182_value; // @[ChiselImProc.scala 346:25]
  reg [1:0] lineBuffer_183_grad_dir; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_183_value; // @[ChiselImProc.scala 346:25]
  reg [1:0] lineBuffer_184_grad_dir; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_184_value; // @[ChiselImProc.scala 346:25]
  reg [1:0] lineBuffer_185_grad_dir; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_185_value; // @[ChiselImProc.scala 346:25]
  reg [1:0] lineBuffer_186_grad_dir; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_186_value; // @[ChiselImProc.scala 346:25]
  reg [1:0] lineBuffer_187_grad_dir; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_187_value; // @[ChiselImProc.scala 346:25]
  reg [1:0] lineBuffer_188_grad_dir; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_188_value; // @[ChiselImProc.scala 346:25]
  reg [1:0] lineBuffer_189_grad_dir; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_189_value; // @[ChiselImProc.scala 346:25]
  reg [1:0] lineBuffer_190_grad_dir; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_190_value; // @[ChiselImProc.scala 346:25]
  reg [1:0] lineBuffer_191_grad_dir; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_191_value; // @[ChiselImProc.scala 346:25]
  reg [1:0] lineBuffer_192_grad_dir; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_192_value; // @[ChiselImProc.scala 346:25]
  reg [1:0] lineBuffer_193_grad_dir; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_193_value; // @[ChiselImProc.scala 346:25]
  reg [1:0] lineBuffer_194_grad_dir; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_194_value; // @[ChiselImProc.scala 346:25]
  reg [1:0] lineBuffer_195_grad_dir; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_195_value; // @[ChiselImProc.scala 346:25]
  reg [1:0] lineBuffer_196_grad_dir; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_196_value; // @[ChiselImProc.scala 346:25]
  reg [1:0] lineBuffer_197_grad_dir; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_197_value; // @[ChiselImProc.scala 346:25]
  reg [1:0] lineBuffer_198_grad_dir; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_198_value; // @[ChiselImProc.scala 346:25]
  reg [1:0] lineBuffer_199_grad_dir; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_199_value; // @[ChiselImProc.scala 346:25]
  reg [1:0] lineBuffer_200_grad_dir; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_200_value; // @[ChiselImProc.scala 346:25]
  reg [1:0] lineBuffer_201_grad_dir; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_201_value; // @[ChiselImProc.scala 346:25]
  reg [1:0] lineBuffer_202_grad_dir; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_202_value; // @[ChiselImProc.scala 346:25]
  reg [1:0] lineBuffer_203_grad_dir; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_203_value; // @[ChiselImProc.scala 346:25]
  reg [1:0] lineBuffer_204_grad_dir; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_204_value; // @[ChiselImProc.scala 346:25]
  reg [1:0] lineBuffer_205_grad_dir; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_205_value; // @[ChiselImProc.scala 346:25]
  reg [1:0] lineBuffer_206_grad_dir; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_206_value; // @[ChiselImProc.scala 346:25]
  reg [1:0] lineBuffer_207_grad_dir; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_207_value; // @[ChiselImProc.scala 346:25]
  reg [1:0] lineBuffer_208_grad_dir; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_208_value; // @[ChiselImProc.scala 346:25]
  reg [1:0] lineBuffer_209_grad_dir; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_209_value; // @[ChiselImProc.scala 346:25]
  reg [1:0] lineBuffer_210_grad_dir; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_210_value; // @[ChiselImProc.scala 346:25]
  reg [1:0] lineBuffer_211_grad_dir; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_211_value; // @[ChiselImProc.scala 346:25]
  reg [1:0] lineBuffer_212_grad_dir; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_212_value; // @[ChiselImProc.scala 346:25]
  reg [1:0] lineBuffer_213_grad_dir; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_213_value; // @[ChiselImProc.scala 346:25]
  reg [1:0] lineBuffer_214_grad_dir; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_214_value; // @[ChiselImProc.scala 346:25]
  reg [1:0] lineBuffer_215_grad_dir; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_215_value; // @[ChiselImProc.scala 346:25]
  reg [1:0] lineBuffer_216_grad_dir; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_216_value; // @[ChiselImProc.scala 346:25]
  reg [1:0] lineBuffer_217_grad_dir; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_217_value; // @[ChiselImProc.scala 346:25]
  reg [1:0] lineBuffer_218_grad_dir; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_218_value; // @[ChiselImProc.scala 346:25]
  reg [1:0] lineBuffer_219_grad_dir; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_219_value; // @[ChiselImProc.scala 346:25]
  reg [1:0] lineBuffer_220_grad_dir; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_220_value; // @[ChiselImProc.scala 346:25]
  reg [1:0] lineBuffer_221_grad_dir; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_221_value; // @[ChiselImProc.scala 346:25]
  reg [1:0] lineBuffer_222_grad_dir; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_222_value; // @[ChiselImProc.scala 346:25]
  reg [1:0] lineBuffer_223_grad_dir; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_223_value; // @[ChiselImProc.scala 346:25]
  reg [1:0] lineBuffer_224_grad_dir; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_224_value; // @[ChiselImProc.scala 346:25]
  reg [1:0] lineBuffer_225_grad_dir; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_225_value; // @[ChiselImProc.scala 346:25]
  reg [1:0] lineBuffer_226_grad_dir; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_226_value; // @[ChiselImProc.scala 346:25]
  reg [1:0] lineBuffer_227_grad_dir; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_227_value; // @[ChiselImProc.scala 346:25]
  reg [1:0] lineBuffer_228_grad_dir; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_228_value; // @[ChiselImProc.scala 346:25]
  reg [1:0] lineBuffer_229_grad_dir; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_229_value; // @[ChiselImProc.scala 346:25]
  reg [1:0] lineBuffer_230_grad_dir; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_230_value; // @[ChiselImProc.scala 346:25]
  reg [1:0] lineBuffer_231_grad_dir; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_231_value; // @[ChiselImProc.scala 346:25]
  reg [1:0] lineBuffer_232_grad_dir; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_232_value; // @[ChiselImProc.scala 346:25]
  reg [1:0] lineBuffer_233_grad_dir; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_233_value; // @[ChiselImProc.scala 346:25]
  reg [1:0] lineBuffer_234_grad_dir; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_234_value; // @[ChiselImProc.scala 346:25]
  reg [1:0] lineBuffer_235_grad_dir; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_235_value; // @[ChiselImProc.scala 346:25]
  reg [1:0] lineBuffer_236_grad_dir; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_236_value; // @[ChiselImProc.scala 346:25]
  reg [1:0] lineBuffer_237_grad_dir; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_237_value; // @[ChiselImProc.scala 346:25]
  reg [1:0] lineBuffer_238_grad_dir; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_238_value; // @[ChiselImProc.scala 346:25]
  reg [1:0] lineBuffer_239_grad_dir; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_239_value; // @[ChiselImProc.scala 346:25]
  reg [1:0] lineBuffer_240_grad_dir; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_240_value; // @[ChiselImProc.scala 346:25]
  reg [1:0] lineBuffer_241_grad_dir; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_241_value; // @[ChiselImProc.scala 346:25]
  reg [1:0] lineBuffer_242_grad_dir; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_242_value; // @[ChiselImProc.scala 346:25]
  reg [1:0] lineBuffer_243_grad_dir; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_243_value; // @[ChiselImProc.scala 346:25]
  reg [1:0] lineBuffer_244_grad_dir; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_244_value; // @[ChiselImProc.scala 346:25]
  reg [1:0] lineBuffer_245_grad_dir; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_245_value; // @[ChiselImProc.scala 346:25]
  reg [1:0] lineBuffer_246_grad_dir; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_246_value; // @[ChiselImProc.scala 346:25]
  reg [1:0] lineBuffer_247_grad_dir; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_247_value; // @[ChiselImProc.scala 346:25]
  reg [1:0] lineBuffer_248_grad_dir; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_248_value; // @[ChiselImProc.scala 346:25]
  reg [1:0] lineBuffer_249_grad_dir; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_249_value; // @[ChiselImProc.scala 346:25]
  reg [1:0] lineBuffer_250_grad_dir; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_250_value; // @[ChiselImProc.scala 346:25]
  reg [1:0] lineBuffer_251_grad_dir; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_251_value; // @[ChiselImProc.scala 346:25]
  reg [1:0] lineBuffer_252_grad_dir; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_252_value; // @[ChiselImProc.scala 346:25]
  reg [1:0] lineBuffer_253_grad_dir; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_253_value; // @[ChiselImProc.scala 346:25]
  reg [1:0] lineBuffer_254_grad_dir; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_254_value; // @[ChiselImProc.scala 346:25]
  reg [1:0] lineBuffer_255_grad_dir; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_255_value; // @[ChiselImProc.scala 346:25]
  reg [1:0] lineBuffer_256_grad_dir; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_256_value; // @[ChiselImProc.scala 346:25]
  reg [1:0] lineBuffer_257_grad_dir; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_257_value; // @[ChiselImProc.scala 346:25]
  reg [1:0] lineBuffer_258_grad_dir; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_258_value; // @[ChiselImProc.scala 346:25]
  reg [1:0] lineBuffer_259_grad_dir; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_259_value; // @[ChiselImProc.scala 346:25]
  reg [1:0] lineBuffer_260_grad_dir; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_260_value; // @[ChiselImProc.scala 346:25]
  reg [1:0] lineBuffer_261_grad_dir; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_261_value; // @[ChiselImProc.scala 346:25]
  reg [1:0] lineBuffer_262_grad_dir; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_262_value; // @[ChiselImProc.scala 346:25]
  reg [1:0] lineBuffer_263_grad_dir; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_263_value; // @[ChiselImProc.scala 346:25]
  reg [1:0] lineBuffer_264_grad_dir; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_264_value; // @[ChiselImProc.scala 346:25]
  reg [1:0] lineBuffer_265_grad_dir; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_265_value; // @[ChiselImProc.scala 346:25]
  reg [1:0] lineBuffer_266_grad_dir; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_266_value; // @[ChiselImProc.scala 346:25]
  reg [1:0] lineBuffer_267_grad_dir; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_267_value; // @[ChiselImProc.scala 346:25]
  reg [1:0] lineBuffer_268_grad_dir; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_268_value; // @[ChiselImProc.scala 346:25]
  reg [1:0] lineBuffer_269_grad_dir; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_269_value; // @[ChiselImProc.scala 346:25]
  reg [1:0] lineBuffer_270_grad_dir; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_270_value; // @[ChiselImProc.scala 346:25]
  reg [1:0] lineBuffer_271_grad_dir; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_271_value; // @[ChiselImProc.scala 346:25]
  reg [1:0] lineBuffer_272_grad_dir; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_272_value; // @[ChiselImProc.scala 346:25]
  reg [1:0] lineBuffer_273_grad_dir; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_273_value; // @[ChiselImProc.scala 346:25]
  reg [1:0] lineBuffer_274_grad_dir; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_274_value; // @[ChiselImProc.scala 346:25]
  reg [1:0] lineBuffer_275_grad_dir; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_275_value; // @[ChiselImProc.scala 346:25]
  reg [1:0] lineBuffer_276_grad_dir; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_276_value; // @[ChiselImProc.scala 346:25]
  reg [1:0] lineBuffer_277_grad_dir; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_277_value; // @[ChiselImProc.scala 346:25]
  reg [1:0] lineBuffer_278_grad_dir; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_278_value; // @[ChiselImProc.scala 346:25]
  reg [1:0] lineBuffer_279_grad_dir; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_279_value; // @[ChiselImProc.scala 346:25]
  reg [1:0] lineBuffer_280_grad_dir; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_280_value; // @[ChiselImProc.scala 346:25]
  reg [1:0] lineBuffer_281_grad_dir; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_281_value; // @[ChiselImProc.scala 346:25]
  reg [1:0] lineBuffer_282_grad_dir; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_282_value; // @[ChiselImProc.scala 346:25]
  reg [1:0] lineBuffer_283_grad_dir; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_283_value; // @[ChiselImProc.scala 346:25]
  reg [1:0] lineBuffer_284_grad_dir; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_284_value; // @[ChiselImProc.scala 346:25]
  reg [1:0] lineBuffer_285_grad_dir; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_285_value; // @[ChiselImProc.scala 346:25]
  reg [1:0] lineBuffer_286_grad_dir; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_286_value; // @[ChiselImProc.scala 346:25]
  reg [1:0] lineBuffer_287_grad_dir; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_287_value; // @[ChiselImProc.scala 346:25]
  reg [1:0] lineBuffer_288_grad_dir; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_288_value; // @[ChiselImProc.scala 346:25]
  reg [1:0] lineBuffer_289_grad_dir; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_289_value; // @[ChiselImProc.scala 346:25]
  reg [1:0] lineBuffer_290_grad_dir; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_290_value; // @[ChiselImProc.scala 346:25]
  reg [1:0] lineBuffer_291_grad_dir; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_291_value; // @[ChiselImProc.scala 346:25]
  reg [1:0] lineBuffer_292_grad_dir; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_292_value; // @[ChiselImProc.scala 346:25]
  reg [1:0] lineBuffer_293_grad_dir; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_293_value; // @[ChiselImProc.scala 346:25]
  reg [1:0] lineBuffer_294_grad_dir; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_294_value; // @[ChiselImProc.scala 346:25]
  reg [1:0] lineBuffer_295_grad_dir; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_295_value; // @[ChiselImProc.scala 346:25]
  reg [1:0] lineBuffer_296_grad_dir; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_296_value; // @[ChiselImProc.scala 346:25]
  reg [1:0] lineBuffer_297_grad_dir; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_297_value; // @[ChiselImProc.scala 346:25]
  reg [1:0] lineBuffer_298_grad_dir; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_298_value; // @[ChiselImProc.scala 346:25]
  reg [1:0] lineBuffer_299_grad_dir; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_299_value; // @[ChiselImProc.scala 346:25]
  reg [1:0] lineBuffer_300_grad_dir; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_300_value; // @[ChiselImProc.scala 346:25]
  reg [1:0] lineBuffer_301_grad_dir; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_301_value; // @[ChiselImProc.scala 346:25]
  reg [1:0] lineBuffer_302_grad_dir; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_302_value; // @[ChiselImProc.scala 346:25]
  reg [1:0] lineBuffer_303_grad_dir; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_303_value; // @[ChiselImProc.scala 346:25]
  reg [1:0] lineBuffer_304_grad_dir; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_304_value; // @[ChiselImProc.scala 346:25]
  reg [1:0] lineBuffer_305_grad_dir; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_305_value; // @[ChiselImProc.scala 346:25]
  reg [1:0] lineBuffer_306_grad_dir; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_306_value; // @[ChiselImProc.scala 346:25]
  reg [1:0] lineBuffer_307_grad_dir; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_307_value; // @[ChiselImProc.scala 346:25]
  reg [1:0] lineBuffer_308_grad_dir; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_308_value; // @[ChiselImProc.scala 346:25]
  reg [1:0] lineBuffer_309_grad_dir; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_309_value; // @[ChiselImProc.scala 346:25]
  reg [1:0] lineBuffer_310_grad_dir; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_310_value; // @[ChiselImProc.scala 346:25]
  reg [1:0] lineBuffer_311_grad_dir; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_311_value; // @[ChiselImProc.scala 346:25]
  reg [1:0] lineBuffer_312_grad_dir; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_312_value; // @[ChiselImProc.scala 346:25]
  reg [1:0] lineBuffer_313_grad_dir; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_313_value; // @[ChiselImProc.scala 346:25]
  reg [1:0] lineBuffer_314_grad_dir; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_314_value; // @[ChiselImProc.scala 346:25]
  reg [1:0] lineBuffer_315_grad_dir; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_315_value; // @[ChiselImProc.scala 346:25]
  reg [1:0] lineBuffer_316_grad_dir; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_316_value; // @[ChiselImProc.scala 346:25]
  reg [1:0] lineBuffer_317_grad_dir; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_317_value; // @[ChiselImProc.scala 346:25]
  reg [1:0] lineBuffer_318_grad_dir; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_318_value; // @[ChiselImProc.scala 346:25]
  reg [1:0] lineBuffer_319_grad_dir; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_319_value; // @[ChiselImProc.scala 346:25]
  reg [1:0] lineBuffer_320_grad_dir; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_320_value; // @[ChiselImProc.scala 346:25]
  reg [1:0] lineBuffer_321_grad_dir; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_321_value; // @[ChiselImProc.scala 346:25]
  reg [1:0] lineBuffer_322_grad_dir; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_322_value; // @[ChiselImProc.scala 346:25]
  reg [1:0] lineBuffer_323_grad_dir; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_323_value; // @[ChiselImProc.scala 346:25]
  reg [1:0] lineBuffer_324_grad_dir; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_324_value; // @[ChiselImProc.scala 346:25]
  reg [1:0] lineBuffer_325_grad_dir; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_325_value; // @[ChiselImProc.scala 346:25]
  reg [1:0] lineBuffer_326_grad_dir; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_326_value; // @[ChiselImProc.scala 346:25]
  reg [1:0] lineBuffer_327_grad_dir; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_327_value; // @[ChiselImProc.scala 346:25]
  reg [1:0] lineBuffer_328_grad_dir; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_328_value; // @[ChiselImProc.scala 346:25]
  reg [1:0] lineBuffer_329_grad_dir; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_329_value; // @[ChiselImProc.scala 346:25]
  reg [1:0] lineBuffer_330_grad_dir; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_330_value; // @[ChiselImProc.scala 346:25]
  reg [1:0] lineBuffer_331_grad_dir; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_331_value; // @[ChiselImProc.scala 346:25]
  reg [1:0] lineBuffer_332_grad_dir; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_332_value; // @[ChiselImProc.scala 346:25]
  reg [1:0] lineBuffer_333_grad_dir; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_333_value; // @[ChiselImProc.scala 346:25]
  reg [1:0] lineBuffer_334_grad_dir; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_334_value; // @[ChiselImProc.scala 346:25]
  reg [1:0] lineBuffer_335_grad_dir; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_335_value; // @[ChiselImProc.scala 346:25]
  reg [1:0] lineBuffer_336_grad_dir; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_336_value; // @[ChiselImProc.scala 346:25]
  reg [1:0] lineBuffer_337_grad_dir; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_337_value; // @[ChiselImProc.scala 346:25]
  reg [1:0] lineBuffer_338_grad_dir; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_338_value; // @[ChiselImProc.scala 346:25]
  reg [1:0] lineBuffer_339_grad_dir; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_339_value; // @[ChiselImProc.scala 346:25]
  reg [1:0] lineBuffer_340_grad_dir; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_340_value; // @[ChiselImProc.scala 346:25]
  reg [1:0] lineBuffer_341_grad_dir; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_341_value; // @[ChiselImProc.scala 346:25]
  reg [1:0] lineBuffer_342_grad_dir; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_342_value; // @[ChiselImProc.scala 346:25]
  reg [1:0] lineBuffer_343_grad_dir; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_343_value; // @[ChiselImProc.scala 346:25]
  reg [1:0] lineBuffer_344_grad_dir; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_344_value; // @[ChiselImProc.scala 346:25]
  reg [1:0] lineBuffer_345_grad_dir; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_345_value; // @[ChiselImProc.scala 346:25]
  reg [1:0] lineBuffer_346_grad_dir; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_346_value; // @[ChiselImProc.scala 346:25]
  reg [1:0] lineBuffer_347_grad_dir; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_347_value; // @[ChiselImProc.scala 346:25]
  reg [1:0] lineBuffer_348_grad_dir; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_348_value; // @[ChiselImProc.scala 346:25]
  reg [1:0] lineBuffer_349_grad_dir; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_349_value; // @[ChiselImProc.scala 346:25]
  reg [1:0] lineBuffer_350_grad_dir; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_350_value; // @[ChiselImProc.scala 346:25]
  reg [1:0] lineBuffer_351_grad_dir; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_351_value; // @[ChiselImProc.scala 346:25]
  reg [1:0] lineBuffer_352_grad_dir; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_352_value; // @[ChiselImProc.scala 346:25]
  reg [1:0] lineBuffer_353_grad_dir; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_353_value; // @[ChiselImProc.scala 346:25]
  reg [1:0] lineBuffer_354_grad_dir; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_354_value; // @[ChiselImProc.scala 346:25]
  reg [1:0] lineBuffer_355_grad_dir; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_355_value; // @[ChiselImProc.scala 346:25]
  reg [1:0] lineBuffer_356_grad_dir; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_356_value; // @[ChiselImProc.scala 346:25]
  reg [1:0] lineBuffer_357_grad_dir; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_357_value; // @[ChiselImProc.scala 346:25]
  reg [1:0] lineBuffer_358_grad_dir; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_358_value; // @[ChiselImProc.scala 346:25]
  reg [1:0] lineBuffer_359_grad_dir; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_359_value; // @[ChiselImProc.scala 346:25]
  reg [1:0] lineBuffer_360_grad_dir; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_360_value; // @[ChiselImProc.scala 346:25]
  reg [1:0] lineBuffer_361_grad_dir; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_361_value; // @[ChiselImProc.scala 346:25]
  reg [1:0] lineBuffer_362_grad_dir; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_362_value; // @[ChiselImProc.scala 346:25]
  reg [1:0] lineBuffer_363_grad_dir; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_363_value; // @[ChiselImProc.scala 346:25]
  reg [1:0] lineBuffer_364_grad_dir; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_364_value; // @[ChiselImProc.scala 346:25]
  reg [1:0] lineBuffer_365_grad_dir; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_365_value; // @[ChiselImProc.scala 346:25]
  reg [1:0] lineBuffer_366_grad_dir; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_366_value; // @[ChiselImProc.scala 346:25]
  reg [1:0] lineBuffer_367_grad_dir; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_367_value; // @[ChiselImProc.scala 346:25]
  reg [1:0] lineBuffer_368_grad_dir; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_368_value; // @[ChiselImProc.scala 346:25]
  reg [1:0] lineBuffer_369_grad_dir; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_369_value; // @[ChiselImProc.scala 346:25]
  reg [1:0] lineBuffer_370_grad_dir; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_370_value; // @[ChiselImProc.scala 346:25]
  reg [1:0] lineBuffer_371_grad_dir; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_371_value; // @[ChiselImProc.scala 346:25]
  reg [1:0] lineBuffer_372_grad_dir; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_372_value; // @[ChiselImProc.scala 346:25]
  reg [1:0] lineBuffer_373_grad_dir; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_373_value; // @[ChiselImProc.scala 346:25]
  reg [1:0] lineBuffer_374_grad_dir; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_374_value; // @[ChiselImProc.scala 346:25]
  reg [1:0] lineBuffer_375_grad_dir; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_375_value; // @[ChiselImProc.scala 346:25]
  reg [1:0] lineBuffer_376_grad_dir; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_376_value; // @[ChiselImProc.scala 346:25]
  reg [1:0] lineBuffer_377_grad_dir; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_377_value; // @[ChiselImProc.scala 346:25]
  reg [1:0] lineBuffer_378_grad_dir; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_378_value; // @[ChiselImProc.scala 346:25]
  reg [1:0] lineBuffer_379_grad_dir; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_379_value; // @[ChiselImProc.scala 346:25]
  reg [1:0] lineBuffer_380_grad_dir; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_380_value; // @[ChiselImProc.scala 346:25]
  reg [1:0] lineBuffer_381_grad_dir; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_381_value; // @[ChiselImProc.scala 346:25]
  reg [1:0] lineBuffer_382_grad_dir; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_382_value; // @[ChiselImProc.scala 346:25]
  reg [1:0] lineBuffer_383_grad_dir; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_383_value; // @[ChiselImProc.scala 346:25]
  reg [1:0] lineBuffer_384_grad_dir; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_384_value; // @[ChiselImProc.scala 346:25]
  reg [1:0] lineBuffer_385_grad_dir; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_385_value; // @[ChiselImProc.scala 346:25]
  reg [1:0] lineBuffer_386_grad_dir; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_386_value; // @[ChiselImProc.scala 346:25]
  reg [1:0] lineBuffer_387_grad_dir; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_387_value; // @[ChiselImProc.scala 346:25]
  reg [1:0] lineBuffer_388_grad_dir; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_388_value; // @[ChiselImProc.scala 346:25]
  reg [1:0] lineBuffer_389_grad_dir; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_389_value; // @[ChiselImProc.scala 346:25]
  reg [1:0] lineBuffer_390_grad_dir; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_390_value; // @[ChiselImProc.scala 346:25]
  reg [1:0] lineBuffer_391_grad_dir; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_391_value; // @[ChiselImProc.scala 346:25]
  reg [1:0] lineBuffer_392_grad_dir; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_392_value; // @[ChiselImProc.scala 346:25]
  reg [1:0] lineBuffer_393_grad_dir; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_393_value; // @[ChiselImProc.scala 346:25]
  reg [1:0] lineBuffer_394_grad_dir; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_394_value; // @[ChiselImProc.scala 346:25]
  reg [1:0] lineBuffer_395_grad_dir; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_395_value; // @[ChiselImProc.scala 346:25]
  reg [1:0] lineBuffer_396_grad_dir; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_396_value; // @[ChiselImProc.scala 346:25]
  reg [1:0] lineBuffer_397_grad_dir; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_397_value; // @[ChiselImProc.scala 346:25]
  reg [1:0] lineBuffer_398_grad_dir; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_398_value; // @[ChiselImProc.scala 346:25]
  reg [1:0] lineBuffer_399_grad_dir; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_399_value; // @[ChiselImProc.scala 346:25]
  reg [1:0] lineBuffer_400_grad_dir; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_400_value; // @[ChiselImProc.scala 346:25]
  reg [1:0] lineBuffer_401_grad_dir; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_401_value; // @[ChiselImProc.scala 346:25]
  reg [1:0] lineBuffer_402_grad_dir; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_402_value; // @[ChiselImProc.scala 346:25]
  reg [1:0] lineBuffer_403_grad_dir; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_403_value; // @[ChiselImProc.scala 346:25]
  reg [1:0] lineBuffer_404_grad_dir; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_404_value; // @[ChiselImProc.scala 346:25]
  reg [1:0] lineBuffer_405_grad_dir; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_405_value; // @[ChiselImProc.scala 346:25]
  reg [1:0] lineBuffer_406_grad_dir; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_406_value; // @[ChiselImProc.scala 346:25]
  reg [1:0] lineBuffer_407_grad_dir; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_407_value; // @[ChiselImProc.scala 346:25]
  reg [1:0] lineBuffer_408_grad_dir; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_408_value; // @[ChiselImProc.scala 346:25]
  reg [1:0] lineBuffer_409_grad_dir; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_409_value; // @[ChiselImProc.scala 346:25]
  reg [1:0] lineBuffer_410_grad_dir; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_410_value; // @[ChiselImProc.scala 346:25]
  reg [1:0] lineBuffer_411_grad_dir; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_411_value; // @[ChiselImProc.scala 346:25]
  reg [1:0] lineBuffer_412_grad_dir; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_412_value; // @[ChiselImProc.scala 346:25]
  reg [1:0] lineBuffer_413_grad_dir; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_413_value; // @[ChiselImProc.scala 346:25]
  reg [1:0] lineBuffer_414_grad_dir; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_414_value; // @[ChiselImProc.scala 346:25]
  reg [1:0] lineBuffer_415_grad_dir; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_415_value; // @[ChiselImProc.scala 346:25]
  reg [1:0] lineBuffer_416_grad_dir; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_416_value; // @[ChiselImProc.scala 346:25]
  reg [1:0] lineBuffer_417_grad_dir; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_417_value; // @[ChiselImProc.scala 346:25]
  reg [1:0] lineBuffer_418_grad_dir; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_418_value; // @[ChiselImProc.scala 346:25]
  reg [1:0] lineBuffer_419_grad_dir; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_419_value; // @[ChiselImProc.scala 346:25]
  reg [1:0] lineBuffer_420_grad_dir; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_420_value; // @[ChiselImProc.scala 346:25]
  reg [1:0] lineBuffer_421_grad_dir; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_421_value; // @[ChiselImProc.scala 346:25]
  reg [1:0] lineBuffer_422_grad_dir; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_422_value; // @[ChiselImProc.scala 346:25]
  reg [1:0] lineBuffer_423_grad_dir; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_423_value; // @[ChiselImProc.scala 346:25]
  reg [1:0] lineBuffer_424_grad_dir; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_424_value; // @[ChiselImProc.scala 346:25]
  reg [1:0] lineBuffer_425_grad_dir; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_425_value; // @[ChiselImProc.scala 346:25]
  reg [1:0] lineBuffer_426_grad_dir; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_426_value; // @[ChiselImProc.scala 346:25]
  reg [1:0] lineBuffer_427_grad_dir; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_427_value; // @[ChiselImProc.scala 346:25]
  reg [1:0] lineBuffer_428_grad_dir; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_428_value; // @[ChiselImProc.scala 346:25]
  reg [1:0] lineBuffer_429_grad_dir; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_429_value; // @[ChiselImProc.scala 346:25]
  reg [1:0] lineBuffer_430_grad_dir; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_430_value; // @[ChiselImProc.scala 346:25]
  reg [1:0] lineBuffer_431_grad_dir; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_431_value; // @[ChiselImProc.scala 346:25]
  reg [1:0] lineBuffer_432_grad_dir; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_432_value; // @[ChiselImProc.scala 346:25]
  reg [1:0] lineBuffer_433_grad_dir; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_433_value; // @[ChiselImProc.scala 346:25]
  reg [1:0] lineBuffer_434_grad_dir; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_434_value; // @[ChiselImProc.scala 346:25]
  reg [1:0] lineBuffer_435_grad_dir; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_435_value; // @[ChiselImProc.scala 346:25]
  reg [1:0] lineBuffer_436_grad_dir; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_436_value; // @[ChiselImProc.scala 346:25]
  reg [1:0] lineBuffer_437_grad_dir; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_437_value; // @[ChiselImProc.scala 346:25]
  reg [1:0] lineBuffer_438_grad_dir; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_438_value; // @[ChiselImProc.scala 346:25]
  reg [1:0] lineBuffer_439_grad_dir; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_439_value; // @[ChiselImProc.scala 346:25]
  reg [1:0] lineBuffer_440_grad_dir; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_440_value; // @[ChiselImProc.scala 346:25]
  reg [1:0] lineBuffer_441_grad_dir; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_441_value; // @[ChiselImProc.scala 346:25]
  reg [1:0] lineBuffer_442_grad_dir; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_442_value; // @[ChiselImProc.scala 346:25]
  reg [1:0] lineBuffer_443_grad_dir; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_443_value; // @[ChiselImProc.scala 346:25]
  reg [1:0] lineBuffer_444_grad_dir; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_444_value; // @[ChiselImProc.scala 346:25]
  reg [1:0] lineBuffer_445_grad_dir; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_445_value; // @[ChiselImProc.scala 346:25]
  reg [1:0] lineBuffer_446_grad_dir; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_446_value; // @[ChiselImProc.scala 346:25]
  reg [1:0] lineBuffer_447_grad_dir; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_447_value; // @[ChiselImProc.scala 346:25]
  reg [1:0] lineBuffer_448_grad_dir; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_448_value; // @[ChiselImProc.scala 346:25]
  reg [1:0] lineBuffer_449_grad_dir; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_449_value; // @[ChiselImProc.scala 346:25]
  reg [1:0] lineBuffer_450_grad_dir; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_450_value; // @[ChiselImProc.scala 346:25]
  reg [1:0] lineBuffer_451_grad_dir; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_451_value; // @[ChiselImProc.scala 346:25]
  reg [1:0] lineBuffer_452_grad_dir; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_452_value; // @[ChiselImProc.scala 346:25]
  reg [1:0] lineBuffer_453_grad_dir; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_453_value; // @[ChiselImProc.scala 346:25]
  reg [1:0] lineBuffer_454_grad_dir; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_454_value; // @[ChiselImProc.scala 346:25]
  reg [1:0] lineBuffer_455_grad_dir; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_455_value; // @[ChiselImProc.scala 346:25]
  reg [1:0] lineBuffer_456_grad_dir; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_456_value; // @[ChiselImProc.scala 346:25]
  reg [1:0] lineBuffer_457_grad_dir; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_457_value; // @[ChiselImProc.scala 346:25]
  reg [1:0] lineBuffer_458_grad_dir; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_458_value; // @[ChiselImProc.scala 346:25]
  reg [1:0] lineBuffer_459_grad_dir; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_459_value; // @[ChiselImProc.scala 346:25]
  reg [1:0] lineBuffer_460_grad_dir; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_460_value; // @[ChiselImProc.scala 346:25]
  reg [1:0] lineBuffer_461_grad_dir; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_461_value; // @[ChiselImProc.scala 346:25]
  reg [1:0] lineBuffer_462_grad_dir; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_462_value; // @[ChiselImProc.scala 346:25]
  reg [1:0] lineBuffer_463_grad_dir; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_463_value; // @[ChiselImProc.scala 346:25]
  reg [1:0] lineBuffer_464_grad_dir; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_464_value; // @[ChiselImProc.scala 346:25]
  reg [1:0] lineBuffer_465_grad_dir; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_465_value; // @[ChiselImProc.scala 346:25]
  reg [1:0] lineBuffer_466_grad_dir; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_466_value; // @[ChiselImProc.scala 346:25]
  reg [1:0] lineBuffer_467_grad_dir; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_467_value; // @[ChiselImProc.scala 346:25]
  reg [1:0] lineBuffer_468_grad_dir; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_468_value; // @[ChiselImProc.scala 346:25]
  reg [1:0] lineBuffer_469_grad_dir; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_469_value; // @[ChiselImProc.scala 346:25]
  reg [1:0] lineBuffer_470_grad_dir; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_470_value; // @[ChiselImProc.scala 346:25]
  reg [1:0] lineBuffer_471_grad_dir; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_471_value; // @[ChiselImProc.scala 346:25]
  reg [1:0] lineBuffer_472_grad_dir; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_472_value; // @[ChiselImProc.scala 346:25]
  reg [1:0] lineBuffer_473_grad_dir; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_473_value; // @[ChiselImProc.scala 346:25]
  reg [1:0] lineBuffer_474_grad_dir; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_474_value; // @[ChiselImProc.scala 346:25]
  reg [1:0] lineBuffer_475_grad_dir; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_475_value; // @[ChiselImProc.scala 346:25]
  reg [1:0] lineBuffer_476_grad_dir; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_476_value; // @[ChiselImProc.scala 346:25]
  reg [1:0] lineBuffer_477_grad_dir; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_477_value; // @[ChiselImProc.scala 346:25]
  reg [1:0] lineBuffer_478_grad_dir; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_478_value; // @[ChiselImProc.scala 346:25]
  reg [1:0] lineBuffer_479_grad_dir; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_479_value; // @[ChiselImProc.scala 346:25]
  reg [1:0] lineBuffer_480_grad_dir; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_480_value; // @[ChiselImProc.scala 346:25]
  reg [1:0] lineBuffer_481_grad_dir; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_481_value; // @[ChiselImProc.scala 346:25]
  reg [1:0] lineBuffer_482_grad_dir; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_482_value; // @[ChiselImProc.scala 346:25]
  reg [1:0] lineBuffer_483_grad_dir; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_483_value; // @[ChiselImProc.scala 346:25]
  reg [1:0] lineBuffer_484_grad_dir; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_484_value; // @[ChiselImProc.scala 346:25]
  reg [1:0] lineBuffer_485_grad_dir; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_485_value; // @[ChiselImProc.scala 346:25]
  reg [1:0] lineBuffer_486_grad_dir; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_486_value; // @[ChiselImProc.scala 346:25]
  reg [1:0] lineBuffer_487_grad_dir; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_487_value; // @[ChiselImProc.scala 346:25]
  reg [1:0] lineBuffer_488_grad_dir; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_488_value; // @[ChiselImProc.scala 346:25]
  reg [1:0] lineBuffer_489_grad_dir; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_489_value; // @[ChiselImProc.scala 346:25]
  reg [1:0] lineBuffer_490_grad_dir; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_490_value; // @[ChiselImProc.scala 346:25]
  reg [1:0] lineBuffer_491_grad_dir; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_491_value; // @[ChiselImProc.scala 346:25]
  reg [1:0] lineBuffer_492_grad_dir; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_492_value; // @[ChiselImProc.scala 346:25]
  reg [1:0] lineBuffer_493_grad_dir; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_493_value; // @[ChiselImProc.scala 346:25]
  reg [1:0] lineBuffer_494_grad_dir; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_494_value; // @[ChiselImProc.scala 346:25]
  reg [1:0] lineBuffer_495_grad_dir; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_495_value; // @[ChiselImProc.scala 346:25]
  reg [1:0] lineBuffer_496_grad_dir; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_496_value; // @[ChiselImProc.scala 346:25]
  reg [1:0] lineBuffer_497_grad_dir; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_497_value; // @[ChiselImProc.scala 346:25]
  reg [1:0] lineBuffer_498_grad_dir; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_498_value; // @[ChiselImProc.scala 346:25]
  reg [1:0] lineBuffer_499_grad_dir; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_499_value; // @[ChiselImProc.scala 346:25]
  reg [1:0] lineBuffer_500_grad_dir; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_500_value; // @[ChiselImProc.scala 346:25]
  reg [1:0] lineBuffer_501_grad_dir; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_501_value; // @[ChiselImProc.scala 346:25]
  reg [1:0] lineBuffer_502_grad_dir; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_502_value; // @[ChiselImProc.scala 346:25]
  reg [1:0] lineBuffer_503_grad_dir; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_503_value; // @[ChiselImProc.scala 346:25]
  reg [1:0] lineBuffer_504_grad_dir; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_504_value; // @[ChiselImProc.scala 346:25]
  reg [1:0] lineBuffer_505_grad_dir; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_505_value; // @[ChiselImProc.scala 346:25]
  reg [1:0] lineBuffer_506_grad_dir; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_506_value; // @[ChiselImProc.scala 346:25]
  reg [1:0] lineBuffer_507_grad_dir; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_507_value; // @[ChiselImProc.scala 346:25]
  reg [1:0] lineBuffer_508_grad_dir; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_508_value; // @[ChiselImProc.scala 346:25]
  reg [1:0] lineBuffer_509_grad_dir; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_509_value; // @[ChiselImProc.scala 346:25]
  reg [1:0] lineBuffer_510_grad_dir; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_510_value; // @[ChiselImProc.scala 346:25]
  reg [1:0] lineBuffer_511_grad_dir; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_511_value; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_512_value; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_513_value; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_514_value; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_515_value; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_516_value; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_517_value; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_518_value; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_519_value; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_520_value; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_521_value; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_522_value; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_523_value; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_524_value; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_525_value; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_526_value; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_527_value; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_528_value; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_529_value; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_530_value; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_531_value; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_532_value; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_533_value; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_534_value; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_535_value; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_536_value; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_537_value; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_538_value; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_539_value; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_540_value; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_541_value; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_542_value; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_543_value; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_544_value; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_545_value; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_546_value; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_547_value; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_548_value; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_549_value; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_550_value; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_551_value; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_552_value; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_553_value; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_554_value; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_555_value; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_556_value; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_557_value; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_558_value; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_559_value; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_560_value; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_561_value; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_562_value; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_563_value; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_564_value; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_565_value; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_566_value; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_567_value; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_568_value; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_569_value; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_570_value; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_571_value; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_572_value; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_573_value; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_574_value; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_575_value; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_576_value; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_577_value; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_578_value; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_579_value; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_580_value; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_581_value; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_582_value; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_583_value; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_584_value; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_585_value; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_586_value; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_587_value; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_588_value; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_589_value; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_590_value; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_591_value; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_592_value; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_593_value; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_594_value; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_595_value; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_596_value; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_597_value; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_598_value; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_599_value; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_600_value; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_601_value; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_602_value; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_603_value; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_604_value; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_605_value; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_606_value; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_607_value; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_608_value; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_609_value; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_610_value; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_611_value; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_612_value; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_613_value; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_614_value; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_615_value; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_616_value; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_617_value; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_618_value; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_619_value; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_620_value; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_621_value; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_622_value; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_623_value; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_624_value; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_625_value; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_626_value; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_627_value; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_628_value; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_629_value; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_630_value; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_631_value; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_632_value; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_633_value; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_634_value; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_635_value; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_636_value; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_637_value; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_638_value; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_639_value; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_640_value; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_641_value; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_642_value; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_643_value; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_644_value; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_645_value; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_646_value; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_647_value; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_648_value; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_649_value; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_650_value; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_651_value; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_652_value; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_653_value; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_654_value; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_655_value; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_656_value; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_657_value; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_658_value; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_659_value; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_660_value; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_661_value; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_662_value; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_663_value; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_664_value; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_665_value; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_666_value; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_667_value; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_668_value; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_669_value; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_670_value; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_671_value; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_672_value; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_673_value; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_674_value; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_675_value; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_676_value; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_677_value; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_678_value; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_679_value; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_680_value; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_681_value; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_682_value; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_683_value; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_684_value; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_685_value; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_686_value; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_687_value; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_688_value; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_689_value; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_690_value; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_691_value; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_692_value; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_693_value; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_694_value; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_695_value; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_696_value; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_697_value; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_698_value; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_699_value; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_700_value; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_701_value; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_702_value; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_703_value; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_704_value; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_705_value; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_706_value; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_707_value; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_708_value; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_709_value; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_710_value; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_711_value; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_712_value; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_713_value; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_714_value; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_715_value; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_716_value; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_717_value; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_718_value; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_719_value; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_720_value; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_721_value; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_722_value; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_723_value; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_724_value; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_725_value; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_726_value; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_727_value; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_728_value; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_729_value; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_730_value; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_731_value; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_732_value; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_733_value; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_734_value; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_735_value; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_736_value; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_737_value; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_738_value; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_739_value; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_740_value; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_741_value; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_742_value; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_743_value; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_744_value; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_745_value; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_746_value; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_747_value; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_748_value; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_749_value; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_750_value; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_751_value; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_752_value; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_753_value; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_754_value; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_755_value; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_756_value; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_757_value; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_758_value; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_759_value; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_760_value; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_761_value; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_762_value; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_763_value; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_764_value; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_765_value; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_766_value; // @[ChiselImProc.scala 346:25]
  reg [7:0] lineBuffer_767_value; // @[ChiselImProc.scala 346:25]
  reg [7:0] windowBuffer_0_value; // @[ChiselImProc.scala 347:27]
  reg [7:0] windowBuffer_1_value; // @[ChiselImProc.scala 347:27]
  reg [7:0] windowBuffer_2_value; // @[ChiselImProc.scala 347:27]
  reg [7:0] windowBuffer_3_value; // @[ChiselImProc.scala 347:27]
  reg [1:0] windowBuffer_4_grad_dir; // @[ChiselImProc.scala 347:27]
  reg [7:0] windowBuffer_4_value; // @[ChiselImProc.scala 347:27]
  reg [1:0] windowBuffer_5_grad_dir; // @[ChiselImProc.scala 347:27]
  reg [7:0] windowBuffer_5_value; // @[ChiselImProc.scala 347:27]
  reg [7:0] windowBuffer_6_value; // @[ChiselImProc.scala 347:27]
  reg [7:0] windowBuffer_7_value; // @[ChiselImProc.scala 347:27]
  reg [7:0] windowBuffer_8_value; // @[ChiselImProc.scala 347:27]
  wire  _T = 2'h0 == stateReg; // @[Conditional.scala 37:30]
  wire  _T_1 = 2'h1 == stateReg; // @[Conditional.scala 37:30]
  wire  _T_2 = ~io_enq_valid; // @[ChiselImProc.scala 84:39]
  wire  _T_3 = io_deq_ready & _T_2; // @[ChiselImProc.scala 84:36]
  wire  _T_4 = io_deq_ready & io_enq_valid; // @[ChiselImProc.scala 87:42]
  wire  _T_5 = ~io_deq_ready; // @[ChiselImProc.scala 92:29]
  wire  _T_6 = _T_5 & io_enq_valid; // @[ChiselImProc.scala 92:43]
  wire  _T_7 = 2'h2 == stateReg; // @[Conditional.scala 37:30]
  wire  _T_8 = 2'h3 == stateReg; // @[Conditional.scala 37:30]
  wire  _T_9 = stateReg == 2'h0; // @[ChiselImProc.scala 116:35]
  wire  _T_10 = stateReg == 2'h1; // @[ChiselImProc.scala 116:57]
  wire  _T_11 = _T_9 | _T_10; // @[ChiselImProc.scala 116:45]
  wire  _T_12 = stateReg == 2'h3; // @[ChiselImProc.scala 116:77]
  wire  _T_15 = stateReg == 2'h2; // @[ChiselImProc.scala 117:55]
  wire  _T_16 = _T_10 | _T_15; // @[ChiselImProc.scala 117:43]
  wire  sel = _T_16 & io_deq_ready; // @[ChiselImProc.scala 352:45]
  wire  _T_798 = 2'h0 == windowBuffer_4_grad_dir; // @[Conditional.scala 37:30]
  wire  _T_799 = windowBuffer_4_value < windowBuffer_3_value; // @[ChiselImProc.scala 373:29]
  wire  _T_800 = windowBuffer_4_value < windowBuffer_5_value; // @[ChiselImProc.scala 373:84]
  wire  _T_801 = _T_799 | _T_800; // @[ChiselImProc.scala 373:71]
  wire [7:0] _GEN_56 = _T_801 ? 8'h0 : windowBuffer_4_value; // @[ChiselImProc.scala 373:127]
  wire  _T_802 = 2'h1 == windowBuffer_4_grad_dir; // @[Conditional.scala 37:30]
  wire  _T_803 = windowBuffer_4_value < windowBuffer_0_value; // @[ChiselImProc.scala 381:28]
  wire  _T_804 = windowBuffer_4_value < windowBuffer_8_value; // @[ChiselImProc.scala 381:65]
  wire  _T_805 = _T_803 | _T_804; // @[ChiselImProc.scala 381:52]
  wire [7:0] _GEN_57 = _T_805 ? 8'h0 : windowBuffer_4_value; // @[ChiselImProc.scala 381:114]
  wire  _T_806 = 2'h2 == windowBuffer_4_grad_dir; // @[Conditional.scala 37:30]
  wire  _T_807 = windowBuffer_4_value < windowBuffer_1_value; // @[ChiselImProc.scala 389:28]
  wire  _T_808 = windowBuffer_4_value < windowBuffer_7_value; // @[ChiselImProc.scala 389:93]
  wire  _T_809 = _T_807 | _T_808; // @[ChiselImProc.scala 389:80]
  wire [7:0] _GEN_58 = _T_809 ? 8'h0 : windowBuffer_4_value; // @[ChiselImProc.scala 389:146]
  wire  _T_810 = 2'h3 == windowBuffer_4_grad_dir; // @[Conditional.scala 37:30]
  wire  _T_811 = windowBuffer_4_value < windowBuffer_2_value; // @[ChiselImProc.scala 397:28]
  wire  _T_812 = windowBuffer_4_value < windowBuffer_6_value; // @[ChiselImProc.scala 397:77]
  wire  _T_813 = _T_811 | _T_812; // @[ChiselImProc.scala 397:64]
  wire [7:0] _GEN_59 = _T_813 ? 8'h0 : windowBuffer_4_value; // @[ChiselImProc.scala 397:128]
  wire [7:0] _GEN_60 = _T_810 ? _GEN_59 : 8'h0; // @[Conditional.scala 39:67]
  wire [7:0] _GEN_61 = _T_806 ? _GEN_58 : _GEN_60; // @[Conditional.scala 39:67]
  wire [7:0] _GEN_62 = _T_802 ? _GEN_57 : _GEN_61; // @[Conditional.scala 39:67]
  assign io_enq_ready = _T_11 | _T_12; // @[ChiselImProc.scala 116:22]
  assign io_deq_valid = _T_10 | _T_15; // @[ChiselImProc.scala 117:22]
  assign io_deq_bits = _T_798 ? _GEN_56 : _GEN_62; // @[ChiselImProc.scala 405:16]
  assign io_deq_user = userReg; // @[ChiselImProc.scala 114:21]
  assign io_deq_last = lastReg; // @[ChiselImProc.scala 113:21]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  stateReg = _RAND_0[1:0];
  _RAND_1 = {1{`RANDOM}};
  dataReg_grad_dir = _RAND_1[1:0];
  _RAND_2 = {1{`RANDOM}};
  dataReg_value = _RAND_2[7:0];
  _RAND_3 = {1{`RANDOM}};
  shadowReg_grad_dir = _RAND_3[1:0];
  _RAND_4 = {1{`RANDOM}};
  shadowReg_value = _RAND_4[7:0];
  _RAND_5 = {1{`RANDOM}};
  userReg = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  shadowUserReg = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  lastReg = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  shadowLastReg = _RAND_8[0:0];
  _RAND_9 = {1{`RANDOM}};
  lineBuffer_0_grad_dir = _RAND_9[1:0];
  _RAND_10 = {1{`RANDOM}};
  lineBuffer_0_value = _RAND_10[7:0];
  _RAND_11 = {1{`RANDOM}};
  lineBuffer_1_grad_dir = _RAND_11[1:0];
  _RAND_12 = {1{`RANDOM}};
  lineBuffer_1_value = _RAND_12[7:0];
  _RAND_13 = {1{`RANDOM}};
  lineBuffer_2_grad_dir = _RAND_13[1:0];
  _RAND_14 = {1{`RANDOM}};
  lineBuffer_2_value = _RAND_14[7:0];
  _RAND_15 = {1{`RANDOM}};
  lineBuffer_3_grad_dir = _RAND_15[1:0];
  _RAND_16 = {1{`RANDOM}};
  lineBuffer_3_value = _RAND_16[7:0];
  _RAND_17 = {1{`RANDOM}};
  lineBuffer_4_grad_dir = _RAND_17[1:0];
  _RAND_18 = {1{`RANDOM}};
  lineBuffer_4_value = _RAND_18[7:0];
  _RAND_19 = {1{`RANDOM}};
  lineBuffer_5_grad_dir = _RAND_19[1:0];
  _RAND_20 = {1{`RANDOM}};
  lineBuffer_5_value = _RAND_20[7:0];
  _RAND_21 = {1{`RANDOM}};
  lineBuffer_6_grad_dir = _RAND_21[1:0];
  _RAND_22 = {1{`RANDOM}};
  lineBuffer_6_value = _RAND_22[7:0];
  _RAND_23 = {1{`RANDOM}};
  lineBuffer_7_grad_dir = _RAND_23[1:0];
  _RAND_24 = {1{`RANDOM}};
  lineBuffer_7_value = _RAND_24[7:0];
  _RAND_25 = {1{`RANDOM}};
  lineBuffer_8_grad_dir = _RAND_25[1:0];
  _RAND_26 = {1{`RANDOM}};
  lineBuffer_8_value = _RAND_26[7:0];
  _RAND_27 = {1{`RANDOM}};
  lineBuffer_9_grad_dir = _RAND_27[1:0];
  _RAND_28 = {1{`RANDOM}};
  lineBuffer_9_value = _RAND_28[7:0];
  _RAND_29 = {1{`RANDOM}};
  lineBuffer_10_grad_dir = _RAND_29[1:0];
  _RAND_30 = {1{`RANDOM}};
  lineBuffer_10_value = _RAND_30[7:0];
  _RAND_31 = {1{`RANDOM}};
  lineBuffer_11_grad_dir = _RAND_31[1:0];
  _RAND_32 = {1{`RANDOM}};
  lineBuffer_11_value = _RAND_32[7:0];
  _RAND_33 = {1{`RANDOM}};
  lineBuffer_12_grad_dir = _RAND_33[1:0];
  _RAND_34 = {1{`RANDOM}};
  lineBuffer_12_value = _RAND_34[7:0];
  _RAND_35 = {1{`RANDOM}};
  lineBuffer_13_grad_dir = _RAND_35[1:0];
  _RAND_36 = {1{`RANDOM}};
  lineBuffer_13_value = _RAND_36[7:0];
  _RAND_37 = {1{`RANDOM}};
  lineBuffer_14_grad_dir = _RAND_37[1:0];
  _RAND_38 = {1{`RANDOM}};
  lineBuffer_14_value = _RAND_38[7:0];
  _RAND_39 = {1{`RANDOM}};
  lineBuffer_15_grad_dir = _RAND_39[1:0];
  _RAND_40 = {1{`RANDOM}};
  lineBuffer_15_value = _RAND_40[7:0];
  _RAND_41 = {1{`RANDOM}};
  lineBuffer_16_grad_dir = _RAND_41[1:0];
  _RAND_42 = {1{`RANDOM}};
  lineBuffer_16_value = _RAND_42[7:0];
  _RAND_43 = {1{`RANDOM}};
  lineBuffer_17_grad_dir = _RAND_43[1:0];
  _RAND_44 = {1{`RANDOM}};
  lineBuffer_17_value = _RAND_44[7:0];
  _RAND_45 = {1{`RANDOM}};
  lineBuffer_18_grad_dir = _RAND_45[1:0];
  _RAND_46 = {1{`RANDOM}};
  lineBuffer_18_value = _RAND_46[7:0];
  _RAND_47 = {1{`RANDOM}};
  lineBuffer_19_grad_dir = _RAND_47[1:0];
  _RAND_48 = {1{`RANDOM}};
  lineBuffer_19_value = _RAND_48[7:0];
  _RAND_49 = {1{`RANDOM}};
  lineBuffer_20_grad_dir = _RAND_49[1:0];
  _RAND_50 = {1{`RANDOM}};
  lineBuffer_20_value = _RAND_50[7:0];
  _RAND_51 = {1{`RANDOM}};
  lineBuffer_21_grad_dir = _RAND_51[1:0];
  _RAND_52 = {1{`RANDOM}};
  lineBuffer_21_value = _RAND_52[7:0];
  _RAND_53 = {1{`RANDOM}};
  lineBuffer_22_grad_dir = _RAND_53[1:0];
  _RAND_54 = {1{`RANDOM}};
  lineBuffer_22_value = _RAND_54[7:0];
  _RAND_55 = {1{`RANDOM}};
  lineBuffer_23_grad_dir = _RAND_55[1:0];
  _RAND_56 = {1{`RANDOM}};
  lineBuffer_23_value = _RAND_56[7:0];
  _RAND_57 = {1{`RANDOM}};
  lineBuffer_24_grad_dir = _RAND_57[1:0];
  _RAND_58 = {1{`RANDOM}};
  lineBuffer_24_value = _RAND_58[7:0];
  _RAND_59 = {1{`RANDOM}};
  lineBuffer_25_grad_dir = _RAND_59[1:0];
  _RAND_60 = {1{`RANDOM}};
  lineBuffer_25_value = _RAND_60[7:0];
  _RAND_61 = {1{`RANDOM}};
  lineBuffer_26_grad_dir = _RAND_61[1:0];
  _RAND_62 = {1{`RANDOM}};
  lineBuffer_26_value = _RAND_62[7:0];
  _RAND_63 = {1{`RANDOM}};
  lineBuffer_27_grad_dir = _RAND_63[1:0];
  _RAND_64 = {1{`RANDOM}};
  lineBuffer_27_value = _RAND_64[7:0];
  _RAND_65 = {1{`RANDOM}};
  lineBuffer_28_grad_dir = _RAND_65[1:0];
  _RAND_66 = {1{`RANDOM}};
  lineBuffer_28_value = _RAND_66[7:0];
  _RAND_67 = {1{`RANDOM}};
  lineBuffer_29_grad_dir = _RAND_67[1:0];
  _RAND_68 = {1{`RANDOM}};
  lineBuffer_29_value = _RAND_68[7:0];
  _RAND_69 = {1{`RANDOM}};
  lineBuffer_30_grad_dir = _RAND_69[1:0];
  _RAND_70 = {1{`RANDOM}};
  lineBuffer_30_value = _RAND_70[7:0];
  _RAND_71 = {1{`RANDOM}};
  lineBuffer_31_grad_dir = _RAND_71[1:0];
  _RAND_72 = {1{`RANDOM}};
  lineBuffer_31_value = _RAND_72[7:0];
  _RAND_73 = {1{`RANDOM}};
  lineBuffer_32_grad_dir = _RAND_73[1:0];
  _RAND_74 = {1{`RANDOM}};
  lineBuffer_32_value = _RAND_74[7:0];
  _RAND_75 = {1{`RANDOM}};
  lineBuffer_33_grad_dir = _RAND_75[1:0];
  _RAND_76 = {1{`RANDOM}};
  lineBuffer_33_value = _RAND_76[7:0];
  _RAND_77 = {1{`RANDOM}};
  lineBuffer_34_grad_dir = _RAND_77[1:0];
  _RAND_78 = {1{`RANDOM}};
  lineBuffer_34_value = _RAND_78[7:0];
  _RAND_79 = {1{`RANDOM}};
  lineBuffer_35_grad_dir = _RAND_79[1:0];
  _RAND_80 = {1{`RANDOM}};
  lineBuffer_35_value = _RAND_80[7:0];
  _RAND_81 = {1{`RANDOM}};
  lineBuffer_36_grad_dir = _RAND_81[1:0];
  _RAND_82 = {1{`RANDOM}};
  lineBuffer_36_value = _RAND_82[7:0];
  _RAND_83 = {1{`RANDOM}};
  lineBuffer_37_grad_dir = _RAND_83[1:0];
  _RAND_84 = {1{`RANDOM}};
  lineBuffer_37_value = _RAND_84[7:0];
  _RAND_85 = {1{`RANDOM}};
  lineBuffer_38_grad_dir = _RAND_85[1:0];
  _RAND_86 = {1{`RANDOM}};
  lineBuffer_38_value = _RAND_86[7:0];
  _RAND_87 = {1{`RANDOM}};
  lineBuffer_39_grad_dir = _RAND_87[1:0];
  _RAND_88 = {1{`RANDOM}};
  lineBuffer_39_value = _RAND_88[7:0];
  _RAND_89 = {1{`RANDOM}};
  lineBuffer_40_grad_dir = _RAND_89[1:0];
  _RAND_90 = {1{`RANDOM}};
  lineBuffer_40_value = _RAND_90[7:0];
  _RAND_91 = {1{`RANDOM}};
  lineBuffer_41_grad_dir = _RAND_91[1:0];
  _RAND_92 = {1{`RANDOM}};
  lineBuffer_41_value = _RAND_92[7:0];
  _RAND_93 = {1{`RANDOM}};
  lineBuffer_42_grad_dir = _RAND_93[1:0];
  _RAND_94 = {1{`RANDOM}};
  lineBuffer_42_value = _RAND_94[7:0];
  _RAND_95 = {1{`RANDOM}};
  lineBuffer_43_grad_dir = _RAND_95[1:0];
  _RAND_96 = {1{`RANDOM}};
  lineBuffer_43_value = _RAND_96[7:0];
  _RAND_97 = {1{`RANDOM}};
  lineBuffer_44_grad_dir = _RAND_97[1:0];
  _RAND_98 = {1{`RANDOM}};
  lineBuffer_44_value = _RAND_98[7:0];
  _RAND_99 = {1{`RANDOM}};
  lineBuffer_45_grad_dir = _RAND_99[1:0];
  _RAND_100 = {1{`RANDOM}};
  lineBuffer_45_value = _RAND_100[7:0];
  _RAND_101 = {1{`RANDOM}};
  lineBuffer_46_grad_dir = _RAND_101[1:0];
  _RAND_102 = {1{`RANDOM}};
  lineBuffer_46_value = _RAND_102[7:0];
  _RAND_103 = {1{`RANDOM}};
  lineBuffer_47_grad_dir = _RAND_103[1:0];
  _RAND_104 = {1{`RANDOM}};
  lineBuffer_47_value = _RAND_104[7:0];
  _RAND_105 = {1{`RANDOM}};
  lineBuffer_48_grad_dir = _RAND_105[1:0];
  _RAND_106 = {1{`RANDOM}};
  lineBuffer_48_value = _RAND_106[7:0];
  _RAND_107 = {1{`RANDOM}};
  lineBuffer_49_grad_dir = _RAND_107[1:0];
  _RAND_108 = {1{`RANDOM}};
  lineBuffer_49_value = _RAND_108[7:0];
  _RAND_109 = {1{`RANDOM}};
  lineBuffer_50_grad_dir = _RAND_109[1:0];
  _RAND_110 = {1{`RANDOM}};
  lineBuffer_50_value = _RAND_110[7:0];
  _RAND_111 = {1{`RANDOM}};
  lineBuffer_51_grad_dir = _RAND_111[1:0];
  _RAND_112 = {1{`RANDOM}};
  lineBuffer_51_value = _RAND_112[7:0];
  _RAND_113 = {1{`RANDOM}};
  lineBuffer_52_grad_dir = _RAND_113[1:0];
  _RAND_114 = {1{`RANDOM}};
  lineBuffer_52_value = _RAND_114[7:0];
  _RAND_115 = {1{`RANDOM}};
  lineBuffer_53_grad_dir = _RAND_115[1:0];
  _RAND_116 = {1{`RANDOM}};
  lineBuffer_53_value = _RAND_116[7:0];
  _RAND_117 = {1{`RANDOM}};
  lineBuffer_54_grad_dir = _RAND_117[1:0];
  _RAND_118 = {1{`RANDOM}};
  lineBuffer_54_value = _RAND_118[7:0];
  _RAND_119 = {1{`RANDOM}};
  lineBuffer_55_grad_dir = _RAND_119[1:0];
  _RAND_120 = {1{`RANDOM}};
  lineBuffer_55_value = _RAND_120[7:0];
  _RAND_121 = {1{`RANDOM}};
  lineBuffer_56_grad_dir = _RAND_121[1:0];
  _RAND_122 = {1{`RANDOM}};
  lineBuffer_56_value = _RAND_122[7:0];
  _RAND_123 = {1{`RANDOM}};
  lineBuffer_57_grad_dir = _RAND_123[1:0];
  _RAND_124 = {1{`RANDOM}};
  lineBuffer_57_value = _RAND_124[7:0];
  _RAND_125 = {1{`RANDOM}};
  lineBuffer_58_grad_dir = _RAND_125[1:0];
  _RAND_126 = {1{`RANDOM}};
  lineBuffer_58_value = _RAND_126[7:0];
  _RAND_127 = {1{`RANDOM}};
  lineBuffer_59_grad_dir = _RAND_127[1:0];
  _RAND_128 = {1{`RANDOM}};
  lineBuffer_59_value = _RAND_128[7:0];
  _RAND_129 = {1{`RANDOM}};
  lineBuffer_60_grad_dir = _RAND_129[1:0];
  _RAND_130 = {1{`RANDOM}};
  lineBuffer_60_value = _RAND_130[7:0];
  _RAND_131 = {1{`RANDOM}};
  lineBuffer_61_grad_dir = _RAND_131[1:0];
  _RAND_132 = {1{`RANDOM}};
  lineBuffer_61_value = _RAND_132[7:0];
  _RAND_133 = {1{`RANDOM}};
  lineBuffer_62_grad_dir = _RAND_133[1:0];
  _RAND_134 = {1{`RANDOM}};
  lineBuffer_62_value = _RAND_134[7:0];
  _RAND_135 = {1{`RANDOM}};
  lineBuffer_63_grad_dir = _RAND_135[1:0];
  _RAND_136 = {1{`RANDOM}};
  lineBuffer_63_value = _RAND_136[7:0];
  _RAND_137 = {1{`RANDOM}};
  lineBuffer_64_grad_dir = _RAND_137[1:0];
  _RAND_138 = {1{`RANDOM}};
  lineBuffer_64_value = _RAND_138[7:0];
  _RAND_139 = {1{`RANDOM}};
  lineBuffer_65_grad_dir = _RAND_139[1:0];
  _RAND_140 = {1{`RANDOM}};
  lineBuffer_65_value = _RAND_140[7:0];
  _RAND_141 = {1{`RANDOM}};
  lineBuffer_66_grad_dir = _RAND_141[1:0];
  _RAND_142 = {1{`RANDOM}};
  lineBuffer_66_value = _RAND_142[7:0];
  _RAND_143 = {1{`RANDOM}};
  lineBuffer_67_grad_dir = _RAND_143[1:0];
  _RAND_144 = {1{`RANDOM}};
  lineBuffer_67_value = _RAND_144[7:0];
  _RAND_145 = {1{`RANDOM}};
  lineBuffer_68_grad_dir = _RAND_145[1:0];
  _RAND_146 = {1{`RANDOM}};
  lineBuffer_68_value = _RAND_146[7:0];
  _RAND_147 = {1{`RANDOM}};
  lineBuffer_69_grad_dir = _RAND_147[1:0];
  _RAND_148 = {1{`RANDOM}};
  lineBuffer_69_value = _RAND_148[7:0];
  _RAND_149 = {1{`RANDOM}};
  lineBuffer_70_grad_dir = _RAND_149[1:0];
  _RAND_150 = {1{`RANDOM}};
  lineBuffer_70_value = _RAND_150[7:0];
  _RAND_151 = {1{`RANDOM}};
  lineBuffer_71_grad_dir = _RAND_151[1:0];
  _RAND_152 = {1{`RANDOM}};
  lineBuffer_71_value = _RAND_152[7:0];
  _RAND_153 = {1{`RANDOM}};
  lineBuffer_72_grad_dir = _RAND_153[1:0];
  _RAND_154 = {1{`RANDOM}};
  lineBuffer_72_value = _RAND_154[7:0];
  _RAND_155 = {1{`RANDOM}};
  lineBuffer_73_grad_dir = _RAND_155[1:0];
  _RAND_156 = {1{`RANDOM}};
  lineBuffer_73_value = _RAND_156[7:0];
  _RAND_157 = {1{`RANDOM}};
  lineBuffer_74_grad_dir = _RAND_157[1:0];
  _RAND_158 = {1{`RANDOM}};
  lineBuffer_74_value = _RAND_158[7:0];
  _RAND_159 = {1{`RANDOM}};
  lineBuffer_75_grad_dir = _RAND_159[1:0];
  _RAND_160 = {1{`RANDOM}};
  lineBuffer_75_value = _RAND_160[7:0];
  _RAND_161 = {1{`RANDOM}};
  lineBuffer_76_grad_dir = _RAND_161[1:0];
  _RAND_162 = {1{`RANDOM}};
  lineBuffer_76_value = _RAND_162[7:0];
  _RAND_163 = {1{`RANDOM}};
  lineBuffer_77_grad_dir = _RAND_163[1:0];
  _RAND_164 = {1{`RANDOM}};
  lineBuffer_77_value = _RAND_164[7:0];
  _RAND_165 = {1{`RANDOM}};
  lineBuffer_78_grad_dir = _RAND_165[1:0];
  _RAND_166 = {1{`RANDOM}};
  lineBuffer_78_value = _RAND_166[7:0];
  _RAND_167 = {1{`RANDOM}};
  lineBuffer_79_grad_dir = _RAND_167[1:0];
  _RAND_168 = {1{`RANDOM}};
  lineBuffer_79_value = _RAND_168[7:0];
  _RAND_169 = {1{`RANDOM}};
  lineBuffer_80_grad_dir = _RAND_169[1:0];
  _RAND_170 = {1{`RANDOM}};
  lineBuffer_80_value = _RAND_170[7:0];
  _RAND_171 = {1{`RANDOM}};
  lineBuffer_81_grad_dir = _RAND_171[1:0];
  _RAND_172 = {1{`RANDOM}};
  lineBuffer_81_value = _RAND_172[7:0];
  _RAND_173 = {1{`RANDOM}};
  lineBuffer_82_grad_dir = _RAND_173[1:0];
  _RAND_174 = {1{`RANDOM}};
  lineBuffer_82_value = _RAND_174[7:0];
  _RAND_175 = {1{`RANDOM}};
  lineBuffer_83_grad_dir = _RAND_175[1:0];
  _RAND_176 = {1{`RANDOM}};
  lineBuffer_83_value = _RAND_176[7:0];
  _RAND_177 = {1{`RANDOM}};
  lineBuffer_84_grad_dir = _RAND_177[1:0];
  _RAND_178 = {1{`RANDOM}};
  lineBuffer_84_value = _RAND_178[7:0];
  _RAND_179 = {1{`RANDOM}};
  lineBuffer_85_grad_dir = _RAND_179[1:0];
  _RAND_180 = {1{`RANDOM}};
  lineBuffer_85_value = _RAND_180[7:0];
  _RAND_181 = {1{`RANDOM}};
  lineBuffer_86_grad_dir = _RAND_181[1:0];
  _RAND_182 = {1{`RANDOM}};
  lineBuffer_86_value = _RAND_182[7:0];
  _RAND_183 = {1{`RANDOM}};
  lineBuffer_87_grad_dir = _RAND_183[1:0];
  _RAND_184 = {1{`RANDOM}};
  lineBuffer_87_value = _RAND_184[7:0];
  _RAND_185 = {1{`RANDOM}};
  lineBuffer_88_grad_dir = _RAND_185[1:0];
  _RAND_186 = {1{`RANDOM}};
  lineBuffer_88_value = _RAND_186[7:0];
  _RAND_187 = {1{`RANDOM}};
  lineBuffer_89_grad_dir = _RAND_187[1:0];
  _RAND_188 = {1{`RANDOM}};
  lineBuffer_89_value = _RAND_188[7:0];
  _RAND_189 = {1{`RANDOM}};
  lineBuffer_90_grad_dir = _RAND_189[1:0];
  _RAND_190 = {1{`RANDOM}};
  lineBuffer_90_value = _RAND_190[7:0];
  _RAND_191 = {1{`RANDOM}};
  lineBuffer_91_grad_dir = _RAND_191[1:0];
  _RAND_192 = {1{`RANDOM}};
  lineBuffer_91_value = _RAND_192[7:0];
  _RAND_193 = {1{`RANDOM}};
  lineBuffer_92_grad_dir = _RAND_193[1:0];
  _RAND_194 = {1{`RANDOM}};
  lineBuffer_92_value = _RAND_194[7:0];
  _RAND_195 = {1{`RANDOM}};
  lineBuffer_93_grad_dir = _RAND_195[1:0];
  _RAND_196 = {1{`RANDOM}};
  lineBuffer_93_value = _RAND_196[7:0];
  _RAND_197 = {1{`RANDOM}};
  lineBuffer_94_grad_dir = _RAND_197[1:0];
  _RAND_198 = {1{`RANDOM}};
  lineBuffer_94_value = _RAND_198[7:0];
  _RAND_199 = {1{`RANDOM}};
  lineBuffer_95_grad_dir = _RAND_199[1:0];
  _RAND_200 = {1{`RANDOM}};
  lineBuffer_95_value = _RAND_200[7:0];
  _RAND_201 = {1{`RANDOM}};
  lineBuffer_96_grad_dir = _RAND_201[1:0];
  _RAND_202 = {1{`RANDOM}};
  lineBuffer_96_value = _RAND_202[7:0];
  _RAND_203 = {1{`RANDOM}};
  lineBuffer_97_grad_dir = _RAND_203[1:0];
  _RAND_204 = {1{`RANDOM}};
  lineBuffer_97_value = _RAND_204[7:0];
  _RAND_205 = {1{`RANDOM}};
  lineBuffer_98_grad_dir = _RAND_205[1:0];
  _RAND_206 = {1{`RANDOM}};
  lineBuffer_98_value = _RAND_206[7:0];
  _RAND_207 = {1{`RANDOM}};
  lineBuffer_99_grad_dir = _RAND_207[1:0];
  _RAND_208 = {1{`RANDOM}};
  lineBuffer_99_value = _RAND_208[7:0];
  _RAND_209 = {1{`RANDOM}};
  lineBuffer_100_grad_dir = _RAND_209[1:0];
  _RAND_210 = {1{`RANDOM}};
  lineBuffer_100_value = _RAND_210[7:0];
  _RAND_211 = {1{`RANDOM}};
  lineBuffer_101_grad_dir = _RAND_211[1:0];
  _RAND_212 = {1{`RANDOM}};
  lineBuffer_101_value = _RAND_212[7:0];
  _RAND_213 = {1{`RANDOM}};
  lineBuffer_102_grad_dir = _RAND_213[1:0];
  _RAND_214 = {1{`RANDOM}};
  lineBuffer_102_value = _RAND_214[7:0];
  _RAND_215 = {1{`RANDOM}};
  lineBuffer_103_grad_dir = _RAND_215[1:0];
  _RAND_216 = {1{`RANDOM}};
  lineBuffer_103_value = _RAND_216[7:0];
  _RAND_217 = {1{`RANDOM}};
  lineBuffer_104_grad_dir = _RAND_217[1:0];
  _RAND_218 = {1{`RANDOM}};
  lineBuffer_104_value = _RAND_218[7:0];
  _RAND_219 = {1{`RANDOM}};
  lineBuffer_105_grad_dir = _RAND_219[1:0];
  _RAND_220 = {1{`RANDOM}};
  lineBuffer_105_value = _RAND_220[7:0];
  _RAND_221 = {1{`RANDOM}};
  lineBuffer_106_grad_dir = _RAND_221[1:0];
  _RAND_222 = {1{`RANDOM}};
  lineBuffer_106_value = _RAND_222[7:0];
  _RAND_223 = {1{`RANDOM}};
  lineBuffer_107_grad_dir = _RAND_223[1:0];
  _RAND_224 = {1{`RANDOM}};
  lineBuffer_107_value = _RAND_224[7:0];
  _RAND_225 = {1{`RANDOM}};
  lineBuffer_108_grad_dir = _RAND_225[1:0];
  _RAND_226 = {1{`RANDOM}};
  lineBuffer_108_value = _RAND_226[7:0];
  _RAND_227 = {1{`RANDOM}};
  lineBuffer_109_grad_dir = _RAND_227[1:0];
  _RAND_228 = {1{`RANDOM}};
  lineBuffer_109_value = _RAND_228[7:0];
  _RAND_229 = {1{`RANDOM}};
  lineBuffer_110_grad_dir = _RAND_229[1:0];
  _RAND_230 = {1{`RANDOM}};
  lineBuffer_110_value = _RAND_230[7:0];
  _RAND_231 = {1{`RANDOM}};
  lineBuffer_111_grad_dir = _RAND_231[1:0];
  _RAND_232 = {1{`RANDOM}};
  lineBuffer_111_value = _RAND_232[7:0];
  _RAND_233 = {1{`RANDOM}};
  lineBuffer_112_grad_dir = _RAND_233[1:0];
  _RAND_234 = {1{`RANDOM}};
  lineBuffer_112_value = _RAND_234[7:0];
  _RAND_235 = {1{`RANDOM}};
  lineBuffer_113_grad_dir = _RAND_235[1:0];
  _RAND_236 = {1{`RANDOM}};
  lineBuffer_113_value = _RAND_236[7:0];
  _RAND_237 = {1{`RANDOM}};
  lineBuffer_114_grad_dir = _RAND_237[1:0];
  _RAND_238 = {1{`RANDOM}};
  lineBuffer_114_value = _RAND_238[7:0];
  _RAND_239 = {1{`RANDOM}};
  lineBuffer_115_grad_dir = _RAND_239[1:0];
  _RAND_240 = {1{`RANDOM}};
  lineBuffer_115_value = _RAND_240[7:0];
  _RAND_241 = {1{`RANDOM}};
  lineBuffer_116_grad_dir = _RAND_241[1:0];
  _RAND_242 = {1{`RANDOM}};
  lineBuffer_116_value = _RAND_242[7:0];
  _RAND_243 = {1{`RANDOM}};
  lineBuffer_117_grad_dir = _RAND_243[1:0];
  _RAND_244 = {1{`RANDOM}};
  lineBuffer_117_value = _RAND_244[7:0];
  _RAND_245 = {1{`RANDOM}};
  lineBuffer_118_grad_dir = _RAND_245[1:0];
  _RAND_246 = {1{`RANDOM}};
  lineBuffer_118_value = _RAND_246[7:0];
  _RAND_247 = {1{`RANDOM}};
  lineBuffer_119_grad_dir = _RAND_247[1:0];
  _RAND_248 = {1{`RANDOM}};
  lineBuffer_119_value = _RAND_248[7:0];
  _RAND_249 = {1{`RANDOM}};
  lineBuffer_120_grad_dir = _RAND_249[1:0];
  _RAND_250 = {1{`RANDOM}};
  lineBuffer_120_value = _RAND_250[7:0];
  _RAND_251 = {1{`RANDOM}};
  lineBuffer_121_grad_dir = _RAND_251[1:0];
  _RAND_252 = {1{`RANDOM}};
  lineBuffer_121_value = _RAND_252[7:0];
  _RAND_253 = {1{`RANDOM}};
  lineBuffer_122_grad_dir = _RAND_253[1:0];
  _RAND_254 = {1{`RANDOM}};
  lineBuffer_122_value = _RAND_254[7:0];
  _RAND_255 = {1{`RANDOM}};
  lineBuffer_123_grad_dir = _RAND_255[1:0];
  _RAND_256 = {1{`RANDOM}};
  lineBuffer_123_value = _RAND_256[7:0];
  _RAND_257 = {1{`RANDOM}};
  lineBuffer_124_grad_dir = _RAND_257[1:0];
  _RAND_258 = {1{`RANDOM}};
  lineBuffer_124_value = _RAND_258[7:0];
  _RAND_259 = {1{`RANDOM}};
  lineBuffer_125_grad_dir = _RAND_259[1:0];
  _RAND_260 = {1{`RANDOM}};
  lineBuffer_125_value = _RAND_260[7:0];
  _RAND_261 = {1{`RANDOM}};
  lineBuffer_126_grad_dir = _RAND_261[1:0];
  _RAND_262 = {1{`RANDOM}};
  lineBuffer_126_value = _RAND_262[7:0];
  _RAND_263 = {1{`RANDOM}};
  lineBuffer_127_grad_dir = _RAND_263[1:0];
  _RAND_264 = {1{`RANDOM}};
  lineBuffer_127_value = _RAND_264[7:0];
  _RAND_265 = {1{`RANDOM}};
  lineBuffer_128_grad_dir = _RAND_265[1:0];
  _RAND_266 = {1{`RANDOM}};
  lineBuffer_128_value = _RAND_266[7:0];
  _RAND_267 = {1{`RANDOM}};
  lineBuffer_129_grad_dir = _RAND_267[1:0];
  _RAND_268 = {1{`RANDOM}};
  lineBuffer_129_value = _RAND_268[7:0];
  _RAND_269 = {1{`RANDOM}};
  lineBuffer_130_grad_dir = _RAND_269[1:0];
  _RAND_270 = {1{`RANDOM}};
  lineBuffer_130_value = _RAND_270[7:0];
  _RAND_271 = {1{`RANDOM}};
  lineBuffer_131_grad_dir = _RAND_271[1:0];
  _RAND_272 = {1{`RANDOM}};
  lineBuffer_131_value = _RAND_272[7:0];
  _RAND_273 = {1{`RANDOM}};
  lineBuffer_132_grad_dir = _RAND_273[1:0];
  _RAND_274 = {1{`RANDOM}};
  lineBuffer_132_value = _RAND_274[7:0];
  _RAND_275 = {1{`RANDOM}};
  lineBuffer_133_grad_dir = _RAND_275[1:0];
  _RAND_276 = {1{`RANDOM}};
  lineBuffer_133_value = _RAND_276[7:0];
  _RAND_277 = {1{`RANDOM}};
  lineBuffer_134_grad_dir = _RAND_277[1:0];
  _RAND_278 = {1{`RANDOM}};
  lineBuffer_134_value = _RAND_278[7:0];
  _RAND_279 = {1{`RANDOM}};
  lineBuffer_135_grad_dir = _RAND_279[1:0];
  _RAND_280 = {1{`RANDOM}};
  lineBuffer_135_value = _RAND_280[7:0];
  _RAND_281 = {1{`RANDOM}};
  lineBuffer_136_grad_dir = _RAND_281[1:0];
  _RAND_282 = {1{`RANDOM}};
  lineBuffer_136_value = _RAND_282[7:0];
  _RAND_283 = {1{`RANDOM}};
  lineBuffer_137_grad_dir = _RAND_283[1:0];
  _RAND_284 = {1{`RANDOM}};
  lineBuffer_137_value = _RAND_284[7:0];
  _RAND_285 = {1{`RANDOM}};
  lineBuffer_138_grad_dir = _RAND_285[1:0];
  _RAND_286 = {1{`RANDOM}};
  lineBuffer_138_value = _RAND_286[7:0];
  _RAND_287 = {1{`RANDOM}};
  lineBuffer_139_grad_dir = _RAND_287[1:0];
  _RAND_288 = {1{`RANDOM}};
  lineBuffer_139_value = _RAND_288[7:0];
  _RAND_289 = {1{`RANDOM}};
  lineBuffer_140_grad_dir = _RAND_289[1:0];
  _RAND_290 = {1{`RANDOM}};
  lineBuffer_140_value = _RAND_290[7:0];
  _RAND_291 = {1{`RANDOM}};
  lineBuffer_141_grad_dir = _RAND_291[1:0];
  _RAND_292 = {1{`RANDOM}};
  lineBuffer_141_value = _RAND_292[7:0];
  _RAND_293 = {1{`RANDOM}};
  lineBuffer_142_grad_dir = _RAND_293[1:0];
  _RAND_294 = {1{`RANDOM}};
  lineBuffer_142_value = _RAND_294[7:0];
  _RAND_295 = {1{`RANDOM}};
  lineBuffer_143_grad_dir = _RAND_295[1:0];
  _RAND_296 = {1{`RANDOM}};
  lineBuffer_143_value = _RAND_296[7:0];
  _RAND_297 = {1{`RANDOM}};
  lineBuffer_144_grad_dir = _RAND_297[1:0];
  _RAND_298 = {1{`RANDOM}};
  lineBuffer_144_value = _RAND_298[7:0];
  _RAND_299 = {1{`RANDOM}};
  lineBuffer_145_grad_dir = _RAND_299[1:0];
  _RAND_300 = {1{`RANDOM}};
  lineBuffer_145_value = _RAND_300[7:0];
  _RAND_301 = {1{`RANDOM}};
  lineBuffer_146_grad_dir = _RAND_301[1:0];
  _RAND_302 = {1{`RANDOM}};
  lineBuffer_146_value = _RAND_302[7:0];
  _RAND_303 = {1{`RANDOM}};
  lineBuffer_147_grad_dir = _RAND_303[1:0];
  _RAND_304 = {1{`RANDOM}};
  lineBuffer_147_value = _RAND_304[7:0];
  _RAND_305 = {1{`RANDOM}};
  lineBuffer_148_grad_dir = _RAND_305[1:0];
  _RAND_306 = {1{`RANDOM}};
  lineBuffer_148_value = _RAND_306[7:0];
  _RAND_307 = {1{`RANDOM}};
  lineBuffer_149_grad_dir = _RAND_307[1:0];
  _RAND_308 = {1{`RANDOM}};
  lineBuffer_149_value = _RAND_308[7:0];
  _RAND_309 = {1{`RANDOM}};
  lineBuffer_150_grad_dir = _RAND_309[1:0];
  _RAND_310 = {1{`RANDOM}};
  lineBuffer_150_value = _RAND_310[7:0];
  _RAND_311 = {1{`RANDOM}};
  lineBuffer_151_grad_dir = _RAND_311[1:0];
  _RAND_312 = {1{`RANDOM}};
  lineBuffer_151_value = _RAND_312[7:0];
  _RAND_313 = {1{`RANDOM}};
  lineBuffer_152_grad_dir = _RAND_313[1:0];
  _RAND_314 = {1{`RANDOM}};
  lineBuffer_152_value = _RAND_314[7:0];
  _RAND_315 = {1{`RANDOM}};
  lineBuffer_153_grad_dir = _RAND_315[1:0];
  _RAND_316 = {1{`RANDOM}};
  lineBuffer_153_value = _RAND_316[7:0];
  _RAND_317 = {1{`RANDOM}};
  lineBuffer_154_grad_dir = _RAND_317[1:0];
  _RAND_318 = {1{`RANDOM}};
  lineBuffer_154_value = _RAND_318[7:0];
  _RAND_319 = {1{`RANDOM}};
  lineBuffer_155_grad_dir = _RAND_319[1:0];
  _RAND_320 = {1{`RANDOM}};
  lineBuffer_155_value = _RAND_320[7:0];
  _RAND_321 = {1{`RANDOM}};
  lineBuffer_156_grad_dir = _RAND_321[1:0];
  _RAND_322 = {1{`RANDOM}};
  lineBuffer_156_value = _RAND_322[7:0];
  _RAND_323 = {1{`RANDOM}};
  lineBuffer_157_grad_dir = _RAND_323[1:0];
  _RAND_324 = {1{`RANDOM}};
  lineBuffer_157_value = _RAND_324[7:0];
  _RAND_325 = {1{`RANDOM}};
  lineBuffer_158_grad_dir = _RAND_325[1:0];
  _RAND_326 = {1{`RANDOM}};
  lineBuffer_158_value = _RAND_326[7:0];
  _RAND_327 = {1{`RANDOM}};
  lineBuffer_159_grad_dir = _RAND_327[1:0];
  _RAND_328 = {1{`RANDOM}};
  lineBuffer_159_value = _RAND_328[7:0];
  _RAND_329 = {1{`RANDOM}};
  lineBuffer_160_grad_dir = _RAND_329[1:0];
  _RAND_330 = {1{`RANDOM}};
  lineBuffer_160_value = _RAND_330[7:0];
  _RAND_331 = {1{`RANDOM}};
  lineBuffer_161_grad_dir = _RAND_331[1:0];
  _RAND_332 = {1{`RANDOM}};
  lineBuffer_161_value = _RAND_332[7:0];
  _RAND_333 = {1{`RANDOM}};
  lineBuffer_162_grad_dir = _RAND_333[1:0];
  _RAND_334 = {1{`RANDOM}};
  lineBuffer_162_value = _RAND_334[7:0];
  _RAND_335 = {1{`RANDOM}};
  lineBuffer_163_grad_dir = _RAND_335[1:0];
  _RAND_336 = {1{`RANDOM}};
  lineBuffer_163_value = _RAND_336[7:0];
  _RAND_337 = {1{`RANDOM}};
  lineBuffer_164_grad_dir = _RAND_337[1:0];
  _RAND_338 = {1{`RANDOM}};
  lineBuffer_164_value = _RAND_338[7:0];
  _RAND_339 = {1{`RANDOM}};
  lineBuffer_165_grad_dir = _RAND_339[1:0];
  _RAND_340 = {1{`RANDOM}};
  lineBuffer_165_value = _RAND_340[7:0];
  _RAND_341 = {1{`RANDOM}};
  lineBuffer_166_grad_dir = _RAND_341[1:0];
  _RAND_342 = {1{`RANDOM}};
  lineBuffer_166_value = _RAND_342[7:0];
  _RAND_343 = {1{`RANDOM}};
  lineBuffer_167_grad_dir = _RAND_343[1:0];
  _RAND_344 = {1{`RANDOM}};
  lineBuffer_167_value = _RAND_344[7:0];
  _RAND_345 = {1{`RANDOM}};
  lineBuffer_168_grad_dir = _RAND_345[1:0];
  _RAND_346 = {1{`RANDOM}};
  lineBuffer_168_value = _RAND_346[7:0];
  _RAND_347 = {1{`RANDOM}};
  lineBuffer_169_grad_dir = _RAND_347[1:0];
  _RAND_348 = {1{`RANDOM}};
  lineBuffer_169_value = _RAND_348[7:0];
  _RAND_349 = {1{`RANDOM}};
  lineBuffer_170_grad_dir = _RAND_349[1:0];
  _RAND_350 = {1{`RANDOM}};
  lineBuffer_170_value = _RAND_350[7:0];
  _RAND_351 = {1{`RANDOM}};
  lineBuffer_171_grad_dir = _RAND_351[1:0];
  _RAND_352 = {1{`RANDOM}};
  lineBuffer_171_value = _RAND_352[7:0];
  _RAND_353 = {1{`RANDOM}};
  lineBuffer_172_grad_dir = _RAND_353[1:0];
  _RAND_354 = {1{`RANDOM}};
  lineBuffer_172_value = _RAND_354[7:0];
  _RAND_355 = {1{`RANDOM}};
  lineBuffer_173_grad_dir = _RAND_355[1:0];
  _RAND_356 = {1{`RANDOM}};
  lineBuffer_173_value = _RAND_356[7:0];
  _RAND_357 = {1{`RANDOM}};
  lineBuffer_174_grad_dir = _RAND_357[1:0];
  _RAND_358 = {1{`RANDOM}};
  lineBuffer_174_value = _RAND_358[7:0];
  _RAND_359 = {1{`RANDOM}};
  lineBuffer_175_grad_dir = _RAND_359[1:0];
  _RAND_360 = {1{`RANDOM}};
  lineBuffer_175_value = _RAND_360[7:0];
  _RAND_361 = {1{`RANDOM}};
  lineBuffer_176_grad_dir = _RAND_361[1:0];
  _RAND_362 = {1{`RANDOM}};
  lineBuffer_176_value = _RAND_362[7:0];
  _RAND_363 = {1{`RANDOM}};
  lineBuffer_177_grad_dir = _RAND_363[1:0];
  _RAND_364 = {1{`RANDOM}};
  lineBuffer_177_value = _RAND_364[7:0];
  _RAND_365 = {1{`RANDOM}};
  lineBuffer_178_grad_dir = _RAND_365[1:0];
  _RAND_366 = {1{`RANDOM}};
  lineBuffer_178_value = _RAND_366[7:0];
  _RAND_367 = {1{`RANDOM}};
  lineBuffer_179_grad_dir = _RAND_367[1:0];
  _RAND_368 = {1{`RANDOM}};
  lineBuffer_179_value = _RAND_368[7:0];
  _RAND_369 = {1{`RANDOM}};
  lineBuffer_180_grad_dir = _RAND_369[1:0];
  _RAND_370 = {1{`RANDOM}};
  lineBuffer_180_value = _RAND_370[7:0];
  _RAND_371 = {1{`RANDOM}};
  lineBuffer_181_grad_dir = _RAND_371[1:0];
  _RAND_372 = {1{`RANDOM}};
  lineBuffer_181_value = _RAND_372[7:0];
  _RAND_373 = {1{`RANDOM}};
  lineBuffer_182_grad_dir = _RAND_373[1:0];
  _RAND_374 = {1{`RANDOM}};
  lineBuffer_182_value = _RAND_374[7:0];
  _RAND_375 = {1{`RANDOM}};
  lineBuffer_183_grad_dir = _RAND_375[1:0];
  _RAND_376 = {1{`RANDOM}};
  lineBuffer_183_value = _RAND_376[7:0];
  _RAND_377 = {1{`RANDOM}};
  lineBuffer_184_grad_dir = _RAND_377[1:0];
  _RAND_378 = {1{`RANDOM}};
  lineBuffer_184_value = _RAND_378[7:0];
  _RAND_379 = {1{`RANDOM}};
  lineBuffer_185_grad_dir = _RAND_379[1:0];
  _RAND_380 = {1{`RANDOM}};
  lineBuffer_185_value = _RAND_380[7:0];
  _RAND_381 = {1{`RANDOM}};
  lineBuffer_186_grad_dir = _RAND_381[1:0];
  _RAND_382 = {1{`RANDOM}};
  lineBuffer_186_value = _RAND_382[7:0];
  _RAND_383 = {1{`RANDOM}};
  lineBuffer_187_grad_dir = _RAND_383[1:0];
  _RAND_384 = {1{`RANDOM}};
  lineBuffer_187_value = _RAND_384[7:0];
  _RAND_385 = {1{`RANDOM}};
  lineBuffer_188_grad_dir = _RAND_385[1:0];
  _RAND_386 = {1{`RANDOM}};
  lineBuffer_188_value = _RAND_386[7:0];
  _RAND_387 = {1{`RANDOM}};
  lineBuffer_189_grad_dir = _RAND_387[1:0];
  _RAND_388 = {1{`RANDOM}};
  lineBuffer_189_value = _RAND_388[7:0];
  _RAND_389 = {1{`RANDOM}};
  lineBuffer_190_grad_dir = _RAND_389[1:0];
  _RAND_390 = {1{`RANDOM}};
  lineBuffer_190_value = _RAND_390[7:0];
  _RAND_391 = {1{`RANDOM}};
  lineBuffer_191_grad_dir = _RAND_391[1:0];
  _RAND_392 = {1{`RANDOM}};
  lineBuffer_191_value = _RAND_392[7:0];
  _RAND_393 = {1{`RANDOM}};
  lineBuffer_192_grad_dir = _RAND_393[1:0];
  _RAND_394 = {1{`RANDOM}};
  lineBuffer_192_value = _RAND_394[7:0];
  _RAND_395 = {1{`RANDOM}};
  lineBuffer_193_grad_dir = _RAND_395[1:0];
  _RAND_396 = {1{`RANDOM}};
  lineBuffer_193_value = _RAND_396[7:0];
  _RAND_397 = {1{`RANDOM}};
  lineBuffer_194_grad_dir = _RAND_397[1:0];
  _RAND_398 = {1{`RANDOM}};
  lineBuffer_194_value = _RAND_398[7:0];
  _RAND_399 = {1{`RANDOM}};
  lineBuffer_195_grad_dir = _RAND_399[1:0];
  _RAND_400 = {1{`RANDOM}};
  lineBuffer_195_value = _RAND_400[7:0];
  _RAND_401 = {1{`RANDOM}};
  lineBuffer_196_grad_dir = _RAND_401[1:0];
  _RAND_402 = {1{`RANDOM}};
  lineBuffer_196_value = _RAND_402[7:0];
  _RAND_403 = {1{`RANDOM}};
  lineBuffer_197_grad_dir = _RAND_403[1:0];
  _RAND_404 = {1{`RANDOM}};
  lineBuffer_197_value = _RAND_404[7:0];
  _RAND_405 = {1{`RANDOM}};
  lineBuffer_198_grad_dir = _RAND_405[1:0];
  _RAND_406 = {1{`RANDOM}};
  lineBuffer_198_value = _RAND_406[7:0];
  _RAND_407 = {1{`RANDOM}};
  lineBuffer_199_grad_dir = _RAND_407[1:0];
  _RAND_408 = {1{`RANDOM}};
  lineBuffer_199_value = _RAND_408[7:0];
  _RAND_409 = {1{`RANDOM}};
  lineBuffer_200_grad_dir = _RAND_409[1:0];
  _RAND_410 = {1{`RANDOM}};
  lineBuffer_200_value = _RAND_410[7:0];
  _RAND_411 = {1{`RANDOM}};
  lineBuffer_201_grad_dir = _RAND_411[1:0];
  _RAND_412 = {1{`RANDOM}};
  lineBuffer_201_value = _RAND_412[7:0];
  _RAND_413 = {1{`RANDOM}};
  lineBuffer_202_grad_dir = _RAND_413[1:0];
  _RAND_414 = {1{`RANDOM}};
  lineBuffer_202_value = _RAND_414[7:0];
  _RAND_415 = {1{`RANDOM}};
  lineBuffer_203_grad_dir = _RAND_415[1:0];
  _RAND_416 = {1{`RANDOM}};
  lineBuffer_203_value = _RAND_416[7:0];
  _RAND_417 = {1{`RANDOM}};
  lineBuffer_204_grad_dir = _RAND_417[1:0];
  _RAND_418 = {1{`RANDOM}};
  lineBuffer_204_value = _RAND_418[7:0];
  _RAND_419 = {1{`RANDOM}};
  lineBuffer_205_grad_dir = _RAND_419[1:0];
  _RAND_420 = {1{`RANDOM}};
  lineBuffer_205_value = _RAND_420[7:0];
  _RAND_421 = {1{`RANDOM}};
  lineBuffer_206_grad_dir = _RAND_421[1:0];
  _RAND_422 = {1{`RANDOM}};
  lineBuffer_206_value = _RAND_422[7:0];
  _RAND_423 = {1{`RANDOM}};
  lineBuffer_207_grad_dir = _RAND_423[1:0];
  _RAND_424 = {1{`RANDOM}};
  lineBuffer_207_value = _RAND_424[7:0];
  _RAND_425 = {1{`RANDOM}};
  lineBuffer_208_grad_dir = _RAND_425[1:0];
  _RAND_426 = {1{`RANDOM}};
  lineBuffer_208_value = _RAND_426[7:0];
  _RAND_427 = {1{`RANDOM}};
  lineBuffer_209_grad_dir = _RAND_427[1:0];
  _RAND_428 = {1{`RANDOM}};
  lineBuffer_209_value = _RAND_428[7:0];
  _RAND_429 = {1{`RANDOM}};
  lineBuffer_210_grad_dir = _RAND_429[1:0];
  _RAND_430 = {1{`RANDOM}};
  lineBuffer_210_value = _RAND_430[7:0];
  _RAND_431 = {1{`RANDOM}};
  lineBuffer_211_grad_dir = _RAND_431[1:0];
  _RAND_432 = {1{`RANDOM}};
  lineBuffer_211_value = _RAND_432[7:0];
  _RAND_433 = {1{`RANDOM}};
  lineBuffer_212_grad_dir = _RAND_433[1:0];
  _RAND_434 = {1{`RANDOM}};
  lineBuffer_212_value = _RAND_434[7:0];
  _RAND_435 = {1{`RANDOM}};
  lineBuffer_213_grad_dir = _RAND_435[1:0];
  _RAND_436 = {1{`RANDOM}};
  lineBuffer_213_value = _RAND_436[7:0];
  _RAND_437 = {1{`RANDOM}};
  lineBuffer_214_grad_dir = _RAND_437[1:0];
  _RAND_438 = {1{`RANDOM}};
  lineBuffer_214_value = _RAND_438[7:0];
  _RAND_439 = {1{`RANDOM}};
  lineBuffer_215_grad_dir = _RAND_439[1:0];
  _RAND_440 = {1{`RANDOM}};
  lineBuffer_215_value = _RAND_440[7:0];
  _RAND_441 = {1{`RANDOM}};
  lineBuffer_216_grad_dir = _RAND_441[1:0];
  _RAND_442 = {1{`RANDOM}};
  lineBuffer_216_value = _RAND_442[7:0];
  _RAND_443 = {1{`RANDOM}};
  lineBuffer_217_grad_dir = _RAND_443[1:0];
  _RAND_444 = {1{`RANDOM}};
  lineBuffer_217_value = _RAND_444[7:0];
  _RAND_445 = {1{`RANDOM}};
  lineBuffer_218_grad_dir = _RAND_445[1:0];
  _RAND_446 = {1{`RANDOM}};
  lineBuffer_218_value = _RAND_446[7:0];
  _RAND_447 = {1{`RANDOM}};
  lineBuffer_219_grad_dir = _RAND_447[1:0];
  _RAND_448 = {1{`RANDOM}};
  lineBuffer_219_value = _RAND_448[7:0];
  _RAND_449 = {1{`RANDOM}};
  lineBuffer_220_grad_dir = _RAND_449[1:0];
  _RAND_450 = {1{`RANDOM}};
  lineBuffer_220_value = _RAND_450[7:0];
  _RAND_451 = {1{`RANDOM}};
  lineBuffer_221_grad_dir = _RAND_451[1:0];
  _RAND_452 = {1{`RANDOM}};
  lineBuffer_221_value = _RAND_452[7:0];
  _RAND_453 = {1{`RANDOM}};
  lineBuffer_222_grad_dir = _RAND_453[1:0];
  _RAND_454 = {1{`RANDOM}};
  lineBuffer_222_value = _RAND_454[7:0];
  _RAND_455 = {1{`RANDOM}};
  lineBuffer_223_grad_dir = _RAND_455[1:0];
  _RAND_456 = {1{`RANDOM}};
  lineBuffer_223_value = _RAND_456[7:0];
  _RAND_457 = {1{`RANDOM}};
  lineBuffer_224_grad_dir = _RAND_457[1:0];
  _RAND_458 = {1{`RANDOM}};
  lineBuffer_224_value = _RAND_458[7:0];
  _RAND_459 = {1{`RANDOM}};
  lineBuffer_225_grad_dir = _RAND_459[1:0];
  _RAND_460 = {1{`RANDOM}};
  lineBuffer_225_value = _RAND_460[7:0];
  _RAND_461 = {1{`RANDOM}};
  lineBuffer_226_grad_dir = _RAND_461[1:0];
  _RAND_462 = {1{`RANDOM}};
  lineBuffer_226_value = _RAND_462[7:0];
  _RAND_463 = {1{`RANDOM}};
  lineBuffer_227_grad_dir = _RAND_463[1:0];
  _RAND_464 = {1{`RANDOM}};
  lineBuffer_227_value = _RAND_464[7:0];
  _RAND_465 = {1{`RANDOM}};
  lineBuffer_228_grad_dir = _RAND_465[1:0];
  _RAND_466 = {1{`RANDOM}};
  lineBuffer_228_value = _RAND_466[7:0];
  _RAND_467 = {1{`RANDOM}};
  lineBuffer_229_grad_dir = _RAND_467[1:0];
  _RAND_468 = {1{`RANDOM}};
  lineBuffer_229_value = _RAND_468[7:0];
  _RAND_469 = {1{`RANDOM}};
  lineBuffer_230_grad_dir = _RAND_469[1:0];
  _RAND_470 = {1{`RANDOM}};
  lineBuffer_230_value = _RAND_470[7:0];
  _RAND_471 = {1{`RANDOM}};
  lineBuffer_231_grad_dir = _RAND_471[1:0];
  _RAND_472 = {1{`RANDOM}};
  lineBuffer_231_value = _RAND_472[7:0];
  _RAND_473 = {1{`RANDOM}};
  lineBuffer_232_grad_dir = _RAND_473[1:0];
  _RAND_474 = {1{`RANDOM}};
  lineBuffer_232_value = _RAND_474[7:0];
  _RAND_475 = {1{`RANDOM}};
  lineBuffer_233_grad_dir = _RAND_475[1:0];
  _RAND_476 = {1{`RANDOM}};
  lineBuffer_233_value = _RAND_476[7:0];
  _RAND_477 = {1{`RANDOM}};
  lineBuffer_234_grad_dir = _RAND_477[1:0];
  _RAND_478 = {1{`RANDOM}};
  lineBuffer_234_value = _RAND_478[7:0];
  _RAND_479 = {1{`RANDOM}};
  lineBuffer_235_grad_dir = _RAND_479[1:0];
  _RAND_480 = {1{`RANDOM}};
  lineBuffer_235_value = _RAND_480[7:0];
  _RAND_481 = {1{`RANDOM}};
  lineBuffer_236_grad_dir = _RAND_481[1:0];
  _RAND_482 = {1{`RANDOM}};
  lineBuffer_236_value = _RAND_482[7:0];
  _RAND_483 = {1{`RANDOM}};
  lineBuffer_237_grad_dir = _RAND_483[1:0];
  _RAND_484 = {1{`RANDOM}};
  lineBuffer_237_value = _RAND_484[7:0];
  _RAND_485 = {1{`RANDOM}};
  lineBuffer_238_grad_dir = _RAND_485[1:0];
  _RAND_486 = {1{`RANDOM}};
  lineBuffer_238_value = _RAND_486[7:0];
  _RAND_487 = {1{`RANDOM}};
  lineBuffer_239_grad_dir = _RAND_487[1:0];
  _RAND_488 = {1{`RANDOM}};
  lineBuffer_239_value = _RAND_488[7:0];
  _RAND_489 = {1{`RANDOM}};
  lineBuffer_240_grad_dir = _RAND_489[1:0];
  _RAND_490 = {1{`RANDOM}};
  lineBuffer_240_value = _RAND_490[7:0];
  _RAND_491 = {1{`RANDOM}};
  lineBuffer_241_grad_dir = _RAND_491[1:0];
  _RAND_492 = {1{`RANDOM}};
  lineBuffer_241_value = _RAND_492[7:0];
  _RAND_493 = {1{`RANDOM}};
  lineBuffer_242_grad_dir = _RAND_493[1:0];
  _RAND_494 = {1{`RANDOM}};
  lineBuffer_242_value = _RAND_494[7:0];
  _RAND_495 = {1{`RANDOM}};
  lineBuffer_243_grad_dir = _RAND_495[1:0];
  _RAND_496 = {1{`RANDOM}};
  lineBuffer_243_value = _RAND_496[7:0];
  _RAND_497 = {1{`RANDOM}};
  lineBuffer_244_grad_dir = _RAND_497[1:0];
  _RAND_498 = {1{`RANDOM}};
  lineBuffer_244_value = _RAND_498[7:0];
  _RAND_499 = {1{`RANDOM}};
  lineBuffer_245_grad_dir = _RAND_499[1:0];
  _RAND_500 = {1{`RANDOM}};
  lineBuffer_245_value = _RAND_500[7:0];
  _RAND_501 = {1{`RANDOM}};
  lineBuffer_246_grad_dir = _RAND_501[1:0];
  _RAND_502 = {1{`RANDOM}};
  lineBuffer_246_value = _RAND_502[7:0];
  _RAND_503 = {1{`RANDOM}};
  lineBuffer_247_grad_dir = _RAND_503[1:0];
  _RAND_504 = {1{`RANDOM}};
  lineBuffer_247_value = _RAND_504[7:0];
  _RAND_505 = {1{`RANDOM}};
  lineBuffer_248_grad_dir = _RAND_505[1:0];
  _RAND_506 = {1{`RANDOM}};
  lineBuffer_248_value = _RAND_506[7:0];
  _RAND_507 = {1{`RANDOM}};
  lineBuffer_249_grad_dir = _RAND_507[1:0];
  _RAND_508 = {1{`RANDOM}};
  lineBuffer_249_value = _RAND_508[7:0];
  _RAND_509 = {1{`RANDOM}};
  lineBuffer_250_grad_dir = _RAND_509[1:0];
  _RAND_510 = {1{`RANDOM}};
  lineBuffer_250_value = _RAND_510[7:0];
  _RAND_511 = {1{`RANDOM}};
  lineBuffer_251_grad_dir = _RAND_511[1:0];
  _RAND_512 = {1{`RANDOM}};
  lineBuffer_251_value = _RAND_512[7:0];
  _RAND_513 = {1{`RANDOM}};
  lineBuffer_252_grad_dir = _RAND_513[1:0];
  _RAND_514 = {1{`RANDOM}};
  lineBuffer_252_value = _RAND_514[7:0];
  _RAND_515 = {1{`RANDOM}};
  lineBuffer_253_grad_dir = _RAND_515[1:0];
  _RAND_516 = {1{`RANDOM}};
  lineBuffer_253_value = _RAND_516[7:0];
  _RAND_517 = {1{`RANDOM}};
  lineBuffer_254_grad_dir = _RAND_517[1:0];
  _RAND_518 = {1{`RANDOM}};
  lineBuffer_254_value = _RAND_518[7:0];
  _RAND_519 = {1{`RANDOM}};
  lineBuffer_255_grad_dir = _RAND_519[1:0];
  _RAND_520 = {1{`RANDOM}};
  lineBuffer_255_value = _RAND_520[7:0];
  _RAND_521 = {1{`RANDOM}};
  lineBuffer_256_grad_dir = _RAND_521[1:0];
  _RAND_522 = {1{`RANDOM}};
  lineBuffer_256_value = _RAND_522[7:0];
  _RAND_523 = {1{`RANDOM}};
  lineBuffer_257_grad_dir = _RAND_523[1:0];
  _RAND_524 = {1{`RANDOM}};
  lineBuffer_257_value = _RAND_524[7:0];
  _RAND_525 = {1{`RANDOM}};
  lineBuffer_258_grad_dir = _RAND_525[1:0];
  _RAND_526 = {1{`RANDOM}};
  lineBuffer_258_value = _RAND_526[7:0];
  _RAND_527 = {1{`RANDOM}};
  lineBuffer_259_grad_dir = _RAND_527[1:0];
  _RAND_528 = {1{`RANDOM}};
  lineBuffer_259_value = _RAND_528[7:0];
  _RAND_529 = {1{`RANDOM}};
  lineBuffer_260_grad_dir = _RAND_529[1:0];
  _RAND_530 = {1{`RANDOM}};
  lineBuffer_260_value = _RAND_530[7:0];
  _RAND_531 = {1{`RANDOM}};
  lineBuffer_261_grad_dir = _RAND_531[1:0];
  _RAND_532 = {1{`RANDOM}};
  lineBuffer_261_value = _RAND_532[7:0];
  _RAND_533 = {1{`RANDOM}};
  lineBuffer_262_grad_dir = _RAND_533[1:0];
  _RAND_534 = {1{`RANDOM}};
  lineBuffer_262_value = _RAND_534[7:0];
  _RAND_535 = {1{`RANDOM}};
  lineBuffer_263_grad_dir = _RAND_535[1:0];
  _RAND_536 = {1{`RANDOM}};
  lineBuffer_263_value = _RAND_536[7:0];
  _RAND_537 = {1{`RANDOM}};
  lineBuffer_264_grad_dir = _RAND_537[1:0];
  _RAND_538 = {1{`RANDOM}};
  lineBuffer_264_value = _RAND_538[7:0];
  _RAND_539 = {1{`RANDOM}};
  lineBuffer_265_grad_dir = _RAND_539[1:0];
  _RAND_540 = {1{`RANDOM}};
  lineBuffer_265_value = _RAND_540[7:0];
  _RAND_541 = {1{`RANDOM}};
  lineBuffer_266_grad_dir = _RAND_541[1:0];
  _RAND_542 = {1{`RANDOM}};
  lineBuffer_266_value = _RAND_542[7:0];
  _RAND_543 = {1{`RANDOM}};
  lineBuffer_267_grad_dir = _RAND_543[1:0];
  _RAND_544 = {1{`RANDOM}};
  lineBuffer_267_value = _RAND_544[7:0];
  _RAND_545 = {1{`RANDOM}};
  lineBuffer_268_grad_dir = _RAND_545[1:0];
  _RAND_546 = {1{`RANDOM}};
  lineBuffer_268_value = _RAND_546[7:0];
  _RAND_547 = {1{`RANDOM}};
  lineBuffer_269_grad_dir = _RAND_547[1:0];
  _RAND_548 = {1{`RANDOM}};
  lineBuffer_269_value = _RAND_548[7:0];
  _RAND_549 = {1{`RANDOM}};
  lineBuffer_270_grad_dir = _RAND_549[1:0];
  _RAND_550 = {1{`RANDOM}};
  lineBuffer_270_value = _RAND_550[7:0];
  _RAND_551 = {1{`RANDOM}};
  lineBuffer_271_grad_dir = _RAND_551[1:0];
  _RAND_552 = {1{`RANDOM}};
  lineBuffer_271_value = _RAND_552[7:0];
  _RAND_553 = {1{`RANDOM}};
  lineBuffer_272_grad_dir = _RAND_553[1:0];
  _RAND_554 = {1{`RANDOM}};
  lineBuffer_272_value = _RAND_554[7:0];
  _RAND_555 = {1{`RANDOM}};
  lineBuffer_273_grad_dir = _RAND_555[1:0];
  _RAND_556 = {1{`RANDOM}};
  lineBuffer_273_value = _RAND_556[7:0];
  _RAND_557 = {1{`RANDOM}};
  lineBuffer_274_grad_dir = _RAND_557[1:0];
  _RAND_558 = {1{`RANDOM}};
  lineBuffer_274_value = _RAND_558[7:0];
  _RAND_559 = {1{`RANDOM}};
  lineBuffer_275_grad_dir = _RAND_559[1:0];
  _RAND_560 = {1{`RANDOM}};
  lineBuffer_275_value = _RAND_560[7:0];
  _RAND_561 = {1{`RANDOM}};
  lineBuffer_276_grad_dir = _RAND_561[1:0];
  _RAND_562 = {1{`RANDOM}};
  lineBuffer_276_value = _RAND_562[7:0];
  _RAND_563 = {1{`RANDOM}};
  lineBuffer_277_grad_dir = _RAND_563[1:0];
  _RAND_564 = {1{`RANDOM}};
  lineBuffer_277_value = _RAND_564[7:0];
  _RAND_565 = {1{`RANDOM}};
  lineBuffer_278_grad_dir = _RAND_565[1:0];
  _RAND_566 = {1{`RANDOM}};
  lineBuffer_278_value = _RAND_566[7:0];
  _RAND_567 = {1{`RANDOM}};
  lineBuffer_279_grad_dir = _RAND_567[1:0];
  _RAND_568 = {1{`RANDOM}};
  lineBuffer_279_value = _RAND_568[7:0];
  _RAND_569 = {1{`RANDOM}};
  lineBuffer_280_grad_dir = _RAND_569[1:0];
  _RAND_570 = {1{`RANDOM}};
  lineBuffer_280_value = _RAND_570[7:0];
  _RAND_571 = {1{`RANDOM}};
  lineBuffer_281_grad_dir = _RAND_571[1:0];
  _RAND_572 = {1{`RANDOM}};
  lineBuffer_281_value = _RAND_572[7:0];
  _RAND_573 = {1{`RANDOM}};
  lineBuffer_282_grad_dir = _RAND_573[1:0];
  _RAND_574 = {1{`RANDOM}};
  lineBuffer_282_value = _RAND_574[7:0];
  _RAND_575 = {1{`RANDOM}};
  lineBuffer_283_grad_dir = _RAND_575[1:0];
  _RAND_576 = {1{`RANDOM}};
  lineBuffer_283_value = _RAND_576[7:0];
  _RAND_577 = {1{`RANDOM}};
  lineBuffer_284_grad_dir = _RAND_577[1:0];
  _RAND_578 = {1{`RANDOM}};
  lineBuffer_284_value = _RAND_578[7:0];
  _RAND_579 = {1{`RANDOM}};
  lineBuffer_285_grad_dir = _RAND_579[1:0];
  _RAND_580 = {1{`RANDOM}};
  lineBuffer_285_value = _RAND_580[7:0];
  _RAND_581 = {1{`RANDOM}};
  lineBuffer_286_grad_dir = _RAND_581[1:0];
  _RAND_582 = {1{`RANDOM}};
  lineBuffer_286_value = _RAND_582[7:0];
  _RAND_583 = {1{`RANDOM}};
  lineBuffer_287_grad_dir = _RAND_583[1:0];
  _RAND_584 = {1{`RANDOM}};
  lineBuffer_287_value = _RAND_584[7:0];
  _RAND_585 = {1{`RANDOM}};
  lineBuffer_288_grad_dir = _RAND_585[1:0];
  _RAND_586 = {1{`RANDOM}};
  lineBuffer_288_value = _RAND_586[7:0];
  _RAND_587 = {1{`RANDOM}};
  lineBuffer_289_grad_dir = _RAND_587[1:0];
  _RAND_588 = {1{`RANDOM}};
  lineBuffer_289_value = _RAND_588[7:0];
  _RAND_589 = {1{`RANDOM}};
  lineBuffer_290_grad_dir = _RAND_589[1:0];
  _RAND_590 = {1{`RANDOM}};
  lineBuffer_290_value = _RAND_590[7:0];
  _RAND_591 = {1{`RANDOM}};
  lineBuffer_291_grad_dir = _RAND_591[1:0];
  _RAND_592 = {1{`RANDOM}};
  lineBuffer_291_value = _RAND_592[7:0];
  _RAND_593 = {1{`RANDOM}};
  lineBuffer_292_grad_dir = _RAND_593[1:0];
  _RAND_594 = {1{`RANDOM}};
  lineBuffer_292_value = _RAND_594[7:0];
  _RAND_595 = {1{`RANDOM}};
  lineBuffer_293_grad_dir = _RAND_595[1:0];
  _RAND_596 = {1{`RANDOM}};
  lineBuffer_293_value = _RAND_596[7:0];
  _RAND_597 = {1{`RANDOM}};
  lineBuffer_294_grad_dir = _RAND_597[1:0];
  _RAND_598 = {1{`RANDOM}};
  lineBuffer_294_value = _RAND_598[7:0];
  _RAND_599 = {1{`RANDOM}};
  lineBuffer_295_grad_dir = _RAND_599[1:0];
  _RAND_600 = {1{`RANDOM}};
  lineBuffer_295_value = _RAND_600[7:0];
  _RAND_601 = {1{`RANDOM}};
  lineBuffer_296_grad_dir = _RAND_601[1:0];
  _RAND_602 = {1{`RANDOM}};
  lineBuffer_296_value = _RAND_602[7:0];
  _RAND_603 = {1{`RANDOM}};
  lineBuffer_297_grad_dir = _RAND_603[1:0];
  _RAND_604 = {1{`RANDOM}};
  lineBuffer_297_value = _RAND_604[7:0];
  _RAND_605 = {1{`RANDOM}};
  lineBuffer_298_grad_dir = _RAND_605[1:0];
  _RAND_606 = {1{`RANDOM}};
  lineBuffer_298_value = _RAND_606[7:0];
  _RAND_607 = {1{`RANDOM}};
  lineBuffer_299_grad_dir = _RAND_607[1:0];
  _RAND_608 = {1{`RANDOM}};
  lineBuffer_299_value = _RAND_608[7:0];
  _RAND_609 = {1{`RANDOM}};
  lineBuffer_300_grad_dir = _RAND_609[1:0];
  _RAND_610 = {1{`RANDOM}};
  lineBuffer_300_value = _RAND_610[7:0];
  _RAND_611 = {1{`RANDOM}};
  lineBuffer_301_grad_dir = _RAND_611[1:0];
  _RAND_612 = {1{`RANDOM}};
  lineBuffer_301_value = _RAND_612[7:0];
  _RAND_613 = {1{`RANDOM}};
  lineBuffer_302_grad_dir = _RAND_613[1:0];
  _RAND_614 = {1{`RANDOM}};
  lineBuffer_302_value = _RAND_614[7:0];
  _RAND_615 = {1{`RANDOM}};
  lineBuffer_303_grad_dir = _RAND_615[1:0];
  _RAND_616 = {1{`RANDOM}};
  lineBuffer_303_value = _RAND_616[7:0];
  _RAND_617 = {1{`RANDOM}};
  lineBuffer_304_grad_dir = _RAND_617[1:0];
  _RAND_618 = {1{`RANDOM}};
  lineBuffer_304_value = _RAND_618[7:0];
  _RAND_619 = {1{`RANDOM}};
  lineBuffer_305_grad_dir = _RAND_619[1:0];
  _RAND_620 = {1{`RANDOM}};
  lineBuffer_305_value = _RAND_620[7:0];
  _RAND_621 = {1{`RANDOM}};
  lineBuffer_306_grad_dir = _RAND_621[1:0];
  _RAND_622 = {1{`RANDOM}};
  lineBuffer_306_value = _RAND_622[7:0];
  _RAND_623 = {1{`RANDOM}};
  lineBuffer_307_grad_dir = _RAND_623[1:0];
  _RAND_624 = {1{`RANDOM}};
  lineBuffer_307_value = _RAND_624[7:0];
  _RAND_625 = {1{`RANDOM}};
  lineBuffer_308_grad_dir = _RAND_625[1:0];
  _RAND_626 = {1{`RANDOM}};
  lineBuffer_308_value = _RAND_626[7:0];
  _RAND_627 = {1{`RANDOM}};
  lineBuffer_309_grad_dir = _RAND_627[1:0];
  _RAND_628 = {1{`RANDOM}};
  lineBuffer_309_value = _RAND_628[7:0];
  _RAND_629 = {1{`RANDOM}};
  lineBuffer_310_grad_dir = _RAND_629[1:0];
  _RAND_630 = {1{`RANDOM}};
  lineBuffer_310_value = _RAND_630[7:0];
  _RAND_631 = {1{`RANDOM}};
  lineBuffer_311_grad_dir = _RAND_631[1:0];
  _RAND_632 = {1{`RANDOM}};
  lineBuffer_311_value = _RAND_632[7:0];
  _RAND_633 = {1{`RANDOM}};
  lineBuffer_312_grad_dir = _RAND_633[1:0];
  _RAND_634 = {1{`RANDOM}};
  lineBuffer_312_value = _RAND_634[7:0];
  _RAND_635 = {1{`RANDOM}};
  lineBuffer_313_grad_dir = _RAND_635[1:0];
  _RAND_636 = {1{`RANDOM}};
  lineBuffer_313_value = _RAND_636[7:0];
  _RAND_637 = {1{`RANDOM}};
  lineBuffer_314_grad_dir = _RAND_637[1:0];
  _RAND_638 = {1{`RANDOM}};
  lineBuffer_314_value = _RAND_638[7:0];
  _RAND_639 = {1{`RANDOM}};
  lineBuffer_315_grad_dir = _RAND_639[1:0];
  _RAND_640 = {1{`RANDOM}};
  lineBuffer_315_value = _RAND_640[7:0];
  _RAND_641 = {1{`RANDOM}};
  lineBuffer_316_grad_dir = _RAND_641[1:0];
  _RAND_642 = {1{`RANDOM}};
  lineBuffer_316_value = _RAND_642[7:0];
  _RAND_643 = {1{`RANDOM}};
  lineBuffer_317_grad_dir = _RAND_643[1:0];
  _RAND_644 = {1{`RANDOM}};
  lineBuffer_317_value = _RAND_644[7:0];
  _RAND_645 = {1{`RANDOM}};
  lineBuffer_318_grad_dir = _RAND_645[1:0];
  _RAND_646 = {1{`RANDOM}};
  lineBuffer_318_value = _RAND_646[7:0];
  _RAND_647 = {1{`RANDOM}};
  lineBuffer_319_grad_dir = _RAND_647[1:0];
  _RAND_648 = {1{`RANDOM}};
  lineBuffer_319_value = _RAND_648[7:0];
  _RAND_649 = {1{`RANDOM}};
  lineBuffer_320_grad_dir = _RAND_649[1:0];
  _RAND_650 = {1{`RANDOM}};
  lineBuffer_320_value = _RAND_650[7:0];
  _RAND_651 = {1{`RANDOM}};
  lineBuffer_321_grad_dir = _RAND_651[1:0];
  _RAND_652 = {1{`RANDOM}};
  lineBuffer_321_value = _RAND_652[7:0];
  _RAND_653 = {1{`RANDOM}};
  lineBuffer_322_grad_dir = _RAND_653[1:0];
  _RAND_654 = {1{`RANDOM}};
  lineBuffer_322_value = _RAND_654[7:0];
  _RAND_655 = {1{`RANDOM}};
  lineBuffer_323_grad_dir = _RAND_655[1:0];
  _RAND_656 = {1{`RANDOM}};
  lineBuffer_323_value = _RAND_656[7:0];
  _RAND_657 = {1{`RANDOM}};
  lineBuffer_324_grad_dir = _RAND_657[1:0];
  _RAND_658 = {1{`RANDOM}};
  lineBuffer_324_value = _RAND_658[7:0];
  _RAND_659 = {1{`RANDOM}};
  lineBuffer_325_grad_dir = _RAND_659[1:0];
  _RAND_660 = {1{`RANDOM}};
  lineBuffer_325_value = _RAND_660[7:0];
  _RAND_661 = {1{`RANDOM}};
  lineBuffer_326_grad_dir = _RAND_661[1:0];
  _RAND_662 = {1{`RANDOM}};
  lineBuffer_326_value = _RAND_662[7:0];
  _RAND_663 = {1{`RANDOM}};
  lineBuffer_327_grad_dir = _RAND_663[1:0];
  _RAND_664 = {1{`RANDOM}};
  lineBuffer_327_value = _RAND_664[7:0];
  _RAND_665 = {1{`RANDOM}};
  lineBuffer_328_grad_dir = _RAND_665[1:0];
  _RAND_666 = {1{`RANDOM}};
  lineBuffer_328_value = _RAND_666[7:0];
  _RAND_667 = {1{`RANDOM}};
  lineBuffer_329_grad_dir = _RAND_667[1:0];
  _RAND_668 = {1{`RANDOM}};
  lineBuffer_329_value = _RAND_668[7:0];
  _RAND_669 = {1{`RANDOM}};
  lineBuffer_330_grad_dir = _RAND_669[1:0];
  _RAND_670 = {1{`RANDOM}};
  lineBuffer_330_value = _RAND_670[7:0];
  _RAND_671 = {1{`RANDOM}};
  lineBuffer_331_grad_dir = _RAND_671[1:0];
  _RAND_672 = {1{`RANDOM}};
  lineBuffer_331_value = _RAND_672[7:0];
  _RAND_673 = {1{`RANDOM}};
  lineBuffer_332_grad_dir = _RAND_673[1:0];
  _RAND_674 = {1{`RANDOM}};
  lineBuffer_332_value = _RAND_674[7:0];
  _RAND_675 = {1{`RANDOM}};
  lineBuffer_333_grad_dir = _RAND_675[1:0];
  _RAND_676 = {1{`RANDOM}};
  lineBuffer_333_value = _RAND_676[7:0];
  _RAND_677 = {1{`RANDOM}};
  lineBuffer_334_grad_dir = _RAND_677[1:0];
  _RAND_678 = {1{`RANDOM}};
  lineBuffer_334_value = _RAND_678[7:0];
  _RAND_679 = {1{`RANDOM}};
  lineBuffer_335_grad_dir = _RAND_679[1:0];
  _RAND_680 = {1{`RANDOM}};
  lineBuffer_335_value = _RAND_680[7:0];
  _RAND_681 = {1{`RANDOM}};
  lineBuffer_336_grad_dir = _RAND_681[1:0];
  _RAND_682 = {1{`RANDOM}};
  lineBuffer_336_value = _RAND_682[7:0];
  _RAND_683 = {1{`RANDOM}};
  lineBuffer_337_grad_dir = _RAND_683[1:0];
  _RAND_684 = {1{`RANDOM}};
  lineBuffer_337_value = _RAND_684[7:0];
  _RAND_685 = {1{`RANDOM}};
  lineBuffer_338_grad_dir = _RAND_685[1:0];
  _RAND_686 = {1{`RANDOM}};
  lineBuffer_338_value = _RAND_686[7:0];
  _RAND_687 = {1{`RANDOM}};
  lineBuffer_339_grad_dir = _RAND_687[1:0];
  _RAND_688 = {1{`RANDOM}};
  lineBuffer_339_value = _RAND_688[7:0];
  _RAND_689 = {1{`RANDOM}};
  lineBuffer_340_grad_dir = _RAND_689[1:0];
  _RAND_690 = {1{`RANDOM}};
  lineBuffer_340_value = _RAND_690[7:0];
  _RAND_691 = {1{`RANDOM}};
  lineBuffer_341_grad_dir = _RAND_691[1:0];
  _RAND_692 = {1{`RANDOM}};
  lineBuffer_341_value = _RAND_692[7:0];
  _RAND_693 = {1{`RANDOM}};
  lineBuffer_342_grad_dir = _RAND_693[1:0];
  _RAND_694 = {1{`RANDOM}};
  lineBuffer_342_value = _RAND_694[7:0];
  _RAND_695 = {1{`RANDOM}};
  lineBuffer_343_grad_dir = _RAND_695[1:0];
  _RAND_696 = {1{`RANDOM}};
  lineBuffer_343_value = _RAND_696[7:0];
  _RAND_697 = {1{`RANDOM}};
  lineBuffer_344_grad_dir = _RAND_697[1:0];
  _RAND_698 = {1{`RANDOM}};
  lineBuffer_344_value = _RAND_698[7:0];
  _RAND_699 = {1{`RANDOM}};
  lineBuffer_345_grad_dir = _RAND_699[1:0];
  _RAND_700 = {1{`RANDOM}};
  lineBuffer_345_value = _RAND_700[7:0];
  _RAND_701 = {1{`RANDOM}};
  lineBuffer_346_grad_dir = _RAND_701[1:0];
  _RAND_702 = {1{`RANDOM}};
  lineBuffer_346_value = _RAND_702[7:0];
  _RAND_703 = {1{`RANDOM}};
  lineBuffer_347_grad_dir = _RAND_703[1:0];
  _RAND_704 = {1{`RANDOM}};
  lineBuffer_347_value = _RAND_704[7:0];
  _RAND_705 = {1{`RANDOM}};
  lineBuffer_348_grad_dir = _RAND_705[1:0];
  _RAND_706 = {1{`RANDOM}};
  lineBuffer_348_value = _RAND_706[7:0];
  _RAND_707 = {1{`RANDOM}};
  lineBuffer_349_grad_dir = _RAND_707[1:0];
  _RAND_708 = {1{`RANDOM}};
  lineBuffer_349_value = _RAND_708[7:0];
  _RAND_709 = {1{`RANDOM}};
  lineBuffer_350_grad_dir = _RAND_709[1:0];
  _RAND_710 = {1{`RANDOM}};
  lineBuffer_350_value = _RAND_710[7:0];
  _RAND_711 = {1{`RANDOM}};
  lineBuffer_351_grad_dir = _RAND_711[1:0];
  _RAND_712 = {1{`RANDOM}};
  lineBuffer_351_value = _RAND_712[7:0];
  _RAND_713 = {1{`RANDOM}};
  lineBuffer_352_grad_dir = _RAND_713[1:0];
  _RAND_714 = {1{`RANDOM}};
  lineBuffer_352_value = _RAND_714[7:0];
  _RAND_715 = {1{`RANDOM}};
  lineBuffer_353_grad_dir = _RAND_715[1:0];
  _RAND_716 = {1{`RANDOM}};
  lineBuffer_353_value = _RAND_716[7:0];
  _RAND_717 = {1{`RANDOM}};
  lineBuffer_354_grad_dir = _RAND_717[1:0];
  _RAND_718 = {1{`RANDOM}};
  lineBuffer_354_value = _RAND_718[7:0];
  _RAND_719 = {1{`RANDOM}};
  lineBuffer_355_grad_dir = _RAND_719[1:0];
  _RAND_720 = {1{`RANDOM}};
  lineBuffer_355_value = _RAND_720[7:0];
  _RAND_721 = {1{`RANDOM}};
  lineBuffer_356_grad_dir = _RAND_721[1:0];
  _RAND_722 = {1{`RANDOM}};
  lineBuffer_356_value = _RAND_722[7:0];
  _RAND_723 = {1{`RANDOM}};
  lineBuffer_357_grad_dir = _RAND_723[1:0];
  _RAND_724 = {1{`RANDOM}};
  lineBuffer_357_value = _RAND_724[7:0];
  _RAND_725 = {1{`RANDOM}};
  lineBuffer_358_grad_dir = _RAND_725[1:0];
  _RAND_726 = {1{`RANDOM}};
  lineBuffer_358_value = _RAND_726[7:0];
  _RAND_727 = {1{`RANDOM}};
  lineBuffer_359_grad_dir = _RAND_727[1:0];
  _RAND_728 = {1{`RANDOM}};
  lineBuffer_359_value = _RAND_728[7:0];
  _RAND_729 = {1{`RANDOM}};
  lineBuffer_360_grad_dir = _RAND_729[1:0];
  _RAND_730 = {1{`RANDOM}};
  lineBuffer_360_value = _RAND_730[7:0];
  _RAND_731 = {1{`RANDOM}};
  lineBuffer_361_grad_dir = _RAND_731[1:0];
  _RAND_732 = {1{`RANDOM}};
  lineBuffer_361_value = _RAND_732[7:0];
  _RAND_733 = {1{`RANDOM}};
  lineBuffer_362_grad_dir = _RAND_733[1:0];
  _RAND_734 = {1{`RANDOM}};
  lineBuffer_362_value = _RAND_734[7:0];
  _RAND_735 = {1{`RANDOM}};
  lineBuffer_363_grad_dir = _RAND_735[1:0];
  _RAND_736 = {1{`RANDOM}};
  lineBuffer_363_value = _RAND_736[7:0];
  _RAND_737 = {1{`RANDOM}};
  lineBuffer_364_grad_dir = _RAND_737[1:0];
  _RAND_738 = {1{`RANDOM}};
  lineBuffer_364_value = _RAND_738[7:0];
  _RAND_739 = {1{`RANDOM}};
  lineBuffer_365_grad_dir = _RAND_739[1:0];
  _RAND_740 = {1{`RANDOM}};
  lineBuffer_365_value = _RAND_740[7:0];
  _RAND_741 = {1{`RANDOM}};
  lineBuffer_366_grad_dir = _RAND_741[1:0];
  _RAND_742 = {1{`RANDOM}};
  lineBuffer_366_value = _RAND_742[7:0];
  _RAND_743 = {1{`RANDOM}};
  lineBuffer_367_grad_dir = _RAND_743[1:0];
  _RAND_744 = {1{`RANDOM}};
  lineBuffer_367_value = _RAND_744[7:0];
  _RAND_745 = {1{`RANDOM}};
  lineBuffer_368_grad_dir = _RAND_745[1:0];
  _RAND_746 = {1{`RANDOM}};
  lineBuffer_368_value = _RAND_746[7:0];
  _RAND_747 = {1{`RANDOM}};
  lineBuffer_369_grad_dir = _RAND_747[1:0];
  _RAND_748 = {1{`RANDOM}};
  lineBuffer_369_value = _RAND_748[7:0];
  _RAND_749 = {1{`RANDOM}};
  lineBuffer_370_grad_dir = _RAND_749[1:0];
  _RAND_750 = {1{`RANDOM}};
  lineBuffer_370_value = _RAND_750[7:0];
  _RAND_751 = {1{`RANDOM}};
  lineBuffer_371_grad_dir = _RAND_751[1:0];
  _RAND_752 = {1{`RANDOM}};
  lineBuffer_371_value = _RAND_752[7:0];
  _RAND_753 = {1{`RANDOM}};
  lineBuffer_372_grad_dir = _RAND_753[1:0];
  _RAND_754 = {1{`RANDOM}};
  lineBuffer_372_value = _RAND_754[7:0];
  _RAND_755 = {1{`RANDOM}};
  lineBuffer_373_grad_dir = _RAND_755[1:0];
  _RAND_756 = {1{`RANDOM}};
  lineBuffer_373_value = _RAND_756[7:0];
  _RAND_757 = {1{`RANDOM}};
  lineBuffer_374_grad_dir = _RAND_757[1:0];
  _RAND_758 = {1{`RANDOM}};
  lineBuffer_374_value = _RAND_758[7:0];
  _RAND_759 = {1{`RANDOM}};
  lineBuffer_375_grad_dir = _RAND_759[1:0];
  _RAND_760 = {1{`RANDOM}};
  lineBuffer_375_value = _RAND_760[7:0];
  _RAND_761 = {1{`RANDOM}};
  lineBuffer_376_grad_dir = _RAND_761[1:0];
  _RAND_762 = {1{`RANDOM}};
  lineBuffer_376_value = _RAND_762[7:0];
  _RAND_763 = {1{`RANDOM}};
  lineBuffer_377_grad_dir = _RAND_763[1:0];
  _RAND_764 = {1{`RANDOM}};
  lineBuffer_377_value = _RAND_764[7:0];
  _RAND_765 = {1{`RANDOM}};
  lineBuffer_378_grad_dir = _RAND_765[1:0];
  _RAND_766 = {1{`RANDOM}};
  lineBuffer_378_value = _RAND_766[7:0];
  _RAND_767 = {1{`RANDOM}};
  lineBuffer_379_grad_dir = _RAND_767[1:0];
  _RAND_768 = {1{`RANDOM}};
  lineBuffer_379_value = _RAND_768[7:0];
  _RAND_769 = {1{`RANDOM}};
  lineBuffer_380_grad_dir = _RAND_769[1:0];
  _RAND_770 = {1{`RANDOM}};
  lineBuffer_380_value = _RAND_770[7:0];
  _RAND_771 = {1{`RANDOM}};
  lineBuffer_381_grad_dir = _RAND_771[1:0];
  _RAND_772 = {1{`RANDOM}};
  lineBuffer_381_value = _RAND_772[7:0];
  _RAND_773 = {1{`RANDOM}};
  lineBuffer_382_grad_dir = _RAND_773[1:0];
  _RAND_774 = {1{`RANDOM}};
  lineBuffer_382_value = _RAND_774[7:0];
  _RAND_775 = {1{`RANDOM}};
  lineBuffer_383_grad_dir = _RAND_775[1:0];
  _RAND_776 = {1{`RANDOM}};
  lineBuffer_383_value = _RAND_776[7:0];
  _RAND_777 = {1{`RANDOM}};
  lineBuffer_384_grad_dir = _RAND_777[1:0];
  _RAND_778 = {1{`RANDOM}};
  lineBuffer_384_value = _RAND_778[7:0];
  _RAND_779 = {1{`RANDOM}};
  lineBuffer_385_grad_dir = _RAND_779[1:0];
  _RAND_780 = {1{`RANDOM}};
  lineBuffer_385_value = _RAND_780[7:0];
  _RAND_781 = {1{`RANDOM}};
  lineBuffer_386_grad_dir = _RAND_781[1:0];
  _RAND_782 = {1{`RANDOM}};
  lineBuffer_386_value = _RAND_782[7:0];
  _RAND_783 = {1{`RANDOM}};
  lineBuffer_387_grad_dir = _RAND_783[1:0];
  _RAND_784 = {1{`RANDOM}};
  lineBuffer_387_value = _RAND_784[7:0];
  _RAND_785 = {1{`RANDOM}};
  lineBuffer_388_grad_dir = _RAND_785[1:0];
  _RAND_786 = {1{`RANDOM}};
  lineBuffer_388_value = _RAND_786[7:0];
  _RAND_787 = {1{`RANDOM}};
  lineBuffer_389_grad_dir = _RAND_787[1:0];
  _RAND_788 = {1{`RANDOM}};
  lineBuffer_389_value = _RAND_788[7:0];
  _RAND_789 = {1{`RANDOM}};
  lineBuffer_390_grad_dir = _RAND_789[1:0];
  _RAND_790 = {1{`RANDOM}};
  lineBuffer_390_value = _RAND_790[7:0];
  _RAND_791 = {1{`RANDOM}};
  lineBuffer_391_grad_dir = _RAND_791[1:0];
  _RAND_792 = {1{`RANDOM}};
  lineBuffer_391_value = _RAND_792[7:0];
  _RAND_793 = {1{`RANDOM}};
  lineBuffer_392_grad_dir = _RAND_793[1:0];
  _RAND_794 = {1{`RANDOM}};
  lineBuffer_392_value = _RAND_794[7:0];
  _RAND_795 = {1{`RANDOM}};
  lineBuffer_393_grad_dir = _RAND_795[1:0];
  _RAND_796 = {1{`RANDOM}};
  lineBuffer_393_value = _RAND_796[7:0];
  _RAND_797 = {1{`RANDOM}};
  lineBuffer_394_grad_dir = _RAND_797[1:0];
  _RAND_798 = {1{`RANDOM}};
  lineBuffer_394_value = _RAND_798[7:0];
  _RAND_799 = {1{`RANDOM}};
  lineBuffer_395_grad_dir = _RAND_799[1:0];
  _RAND_800 = {1{`RANDOM}};
  lineBuffer_395_value = _RAND_800[7:0];
  _RAND_801 = {1{`RANDOM}};
  lineBuffer_396_grad_dir = _RAND_801[1:0];
  _RAND_802 = {1{`RANDOM}};
  lineBuffer_396_value = _RAND_802[7:0];
  _RAND_803 = {1{`RANDOM}};
  lineBuffer_397_grad_dir = _RAND_803[1:0];
  _RAND_804 = {1{`RANDOM}};
  lineBuffer_397_value = _RAND_804[7:0];
  _RAND_805 = {1{`RANDOM}};
  lineBuffer_398_grad_dir = _RAND_805[1:0];
  _RAND_806 = {1{`RANDOM}};
  lineBuffer_398_value = _RAND_806[7:0];
  _RAND_807 = {1{`RANDOM}};
  lineBuffer_399_grad_dir = _RAND_807[1:0];
  _RAND_808 = {1{`RANDOM}};
  lineBuffer_399_value = _RAND_808[7:0];
  _RAND_809 = {1{`RANDOM}};
  lineBuffer_400_grad_dir = _RAND_809[1:0];
  _RAND_810 = {1{`RANDOM}};
  lineBuffer_400_value = _RAND_810[7:0];
  _RAND_811 = {1{`RANDOM}};
  lineBuffer_401_grad_dir = _RAND_811[1:0];
  _RAND_812 = {1{`RANDOM}};
  lineBuffer_401_value = _RAND_812[7:0];
  _RAND_813 = {1{`RANDOM}};
  lineBuffer_402_grad_dir = _RAND_813[1:0];
  _RAND_814 = {1{`RANDOM}};
  lineBuffer_402_value = _RAND_814[7:0];
  _RAND_815 = {1{`RANDOM}};
  lineBuffer_403_grad_dir = _RAND_815[1:0];
  _RAND_816 = {1{`RANDOM}};
  lineBuffer_403_value = _RAND_816[7:0];
  _RAND_817 = {1{`RANDOM}};
  lineBuffer_404_grad_dir = _RAND_817[1:0];
  _RAND_818 = {1{`RANDOM}};
  lineBuffer_404_value = _RAND_818[7:0];
  _RAND_819 = {1{`RANDOM}};
  lineBuffer_405_grad_dir = _RAND_819[1:0];
  _RAND_820 = {1{`RANDOM}};
  lineBuffer_405_value = _RAND_820[7:0];
  _RAND_821 = {1{`RANDOM}};
  lineBuffer_406_grad_dir = _RAND_821[1:0];
  _RAND_822 = {1{`RANDOM}};
  lineBuffer_406_value = _RAND_822[7:0];
  _RAND_823 = {1{`RANDOM}};
  lineBuffer_407_grad_dir = _RAND_823[1:0];
  _RAND_824 = {1{`RANDOM}};
  lineBuffer_407_value = _RAND_824[7:0];
  _RAND_825 = {1{`RANDOM}};
  lineBuffer_408_grad_dir = _RAND_825[1:0];
  _RAND_826 = {1{`RANDOM}};
  lineBuffer_408_value = _RAND_826[7:0];
  _RAND_827 = {1{`RANDOM}};
  lineBuffer_409_grad_dir = _RAND_827[1:0];
  _RAND_828 = {1{`RANDOM}};
  lineBuffer_409_value = _RAND_828[7:0];
  _RAND_829 = {1{`RANDOM}};
  lineBuffer_410_grad_dir = _RAND_829[1:0];
  _RAND_830 = {1{`RANDOM}};
  lineBuffer_410_value = _RAND_830[7:0];
  _RAND_831 = {1{`RANDOM}};
  lineBuffer_411_grad_dir = _RAND_831[1:0];
  _RAND_832 = {1{`RANDOM}};
  lineBuffer_411_value = _RAND_832[7:0];
  _RAND_833 = {1{`RANDOM}};
  lineBuffer_412_grad_dir = _RAND_833[1:0];
  _RAND_834 = {1{`RANDOM}};
  lineBuffer_412_value = _RAND_834[7:0];
  _RAND_835 = {1{`RANDOM}};
  lineBuffer_413_grad_dir = _RAND_835[1:0];
  _RAND_836 = {1{`RANDOM}};
  lineBuffer_413_value = _RAND_836[7:0];
  _RAND_837 = {1{`RANDOM}};
  lineBuffer_414_grad_dir = _RAND_837[1:0];
  _RAND_838 = {1{`RANDOM}};
  lineBuffer_414_value = _RAND_838[7:0];
  _RAND_839 = {1{`RANDOM}};
  lineBuffer_415_grad_dir = _RAND_839[1:0];
  _RAND_840 = {1{`RANDOM}};
  lineBuffer_415_value = _RAND_840[7:0];
  _RAND_841 = {1{`RANDOM}};
  lineBuffer_416_grad_dir = _RAND_841[1:0];
  _RAND_842 = {1{`RANDOM}};
  lineBuffer_416_value = _RAND_842[7:0];
  _RAND_843 = {1{`RANDOM}};
  lineBuffer_417_grad_dir = _RAND_843[1:0];
  _RAND_844 = {1{`RANDOM}};
  lineBuffer_417_value = _RAND_844[7:0];
  _RAND_845 = {1{`RANDOM}};
  lineBuffer_418_grad_dir = _RAND_845[1:0];
  _RAND_846 = {1{`RANDOM}};
  lineBuffer_418_value = _RAND_846[7:0];
  _RAND_847 = {1{`RANDOM}};
  lineBuffer_419_grad_dir = _RAND_847[1:0];
  _RAND_848 = {1{`RANDOM}};
  lineBuffer_419_value = _RAND_848[7:0];
  _RAND_849 = {1{`RANDOM}};
  lineBuffer_420_grad_dir = _RAND_849[1:0];
  _RAND_850 = {1{`RANDOM}};
  lineBuffer_420_value = _RAND_850[7:0];
  _RAND_851 = {1{`RANDOM}};
  lineBuffer_421_grad_dir = _RAND_851[1:0];
  _RAND_852 = {1{`RANDOM}};
  lineBuffer_421_value = _RAND_852[7:0];
  _RAND_853 = {1{`RANDOM}};
  lineBuffer_422_grad_dir = _RAND_853[1:0];
  _RAND_854 = {1{`RANDOM}};
  lineBuffer_422_value = _RAND_854[7:0];
  _RAND_855 = {1{`RANDOM}};
  lineBuffer_423_grad_dir = _RAND_855[1:0];
  _RAND_856 = {1{`RANDOM}};
  lineBuffer_423_value = _RAND_856[7:0];
  _RAND_857 = {1{`RANDOM}};
  lineBuffer_424_grad_dir = _RAND_857[1:0];
  _RAND_858 = {1{`RANDOM}};
  lineBuffer_424_value = _RAND_858[7:0];
  _RAND_859 = {1{`RANDOM}};
  lineBuffer_425_grad_dir = _RAND_859[1:0];
  _RAND_860 = {1{`RANDOM}};
  lineBuffer_425_value = _RAND_860[7:0];
  _RAND_861 = {1{`RANDOM}};
  lineBuffer_426_grad_dir = _RAND_861[1:0];
  _RAND_862 = {1{`RANDOM}};
  lineBuffer_426_value = _RAND_862[7:0];
  _RAND_863 = {1{`RANDOM}};
  lineBuffer_427_grad_dir = _RAND_863[1:0];
  _RAND_864 = {1{`RANDOM}};
  lineBuffer_427_value = _RAND_864[7:0];
  _RAND_865 = {1{`RANDOM}};
  lineBuffer_428_grad_dir = _RAND_865[1:0];
  _RAND_866 = {1{`RANDOM}};
  lineBuffer_428_value = _RAND_866[7:0];
  _RAND_867 = {1{`RANDOM}};
  lineBuffer_429_grad_dir = _RAND_867[1:0];
  _RAND_868 = {1{`RANDOM}};
  lineBuffer_429_value = _RAND_868[7:0];
  _RAND_869 = {1{`RANDOM}};
  lineBuffer_430_grad_dir = _RAND_869[1:0];
  _RAND_870 = {1{`RANDOM}};
  lineBuffer_430_value = _RAND_870[7:0];
  _RAND_871 = {1{`RANDOM}};
  lineBuffer_431_grad_dir = _RAND_871[1:0];
  _RAND_872 = {1{`RANDOM}};
  lineBuffer_431_value = _RAND_872[7:0];
  _RAND_873 = {1{`RANDOM}};
  lineBuffer_432_grad_dir = _RAND_873[1:0];
  _RAND_874 = {1{`RANDOM}};
  lineBuffer_432_value = _RAND_874[7:0];
  _RAND_875 = {1{`RANDOM}};
  lineBuffer_433_grad_dir = _RAND_875[1:0];
  _RAND_876 = {1{`RANDOM}};
  lineBuffer_433_value = _RAND_876[7:0];
  _RAND_877 = {1{`RANDOM}};
  lineBuffer_434_grad_dir = _RAND_877[1:0];
  _RAND_878 = {1{`RANDOM}};
  lineBuffer_434_value = _RAND_878[7:0];
  _RAND_879 = {1{`RANDOM}};
  lineBuffer_435_grad_dir = _RAND_879[1:0];
  _RAND_880 = {1{`RANDOM}};
  lineBuffer_435_value = _RAND_880[7:0];
  _RAND_881 = {1{`RANDOM}};
  lineBuffer_436_grad_dir = _RAND_881[1:0];
  _RAND_882 = {1{`RANDOM}};
  lineBuffer_436_value = _RAND_882[7:0];
  _RAND_883 = {1{`RANDOM}};
  lineBuffer_437_grad_dir = _RAND_883[1:0];
  _RAND_884 = {1{`RANDOM}};
  lineBuffer_437_value = _RAND_884[7:0];
  _RAND_885 = {1{`RANDOM}};
  lineBuffer_438_grad_dir = _RAND_885[1:0];
  _RAND_886 = {1{`RANDOM}};
  lineBuffer_438_value = _RAND_886[7:0];
  _RAND_887 = {1{`RANDOM}};
  lineBuffer_439_grad_dir = _RAND_887[1:0];
  _RAND_888 = {1{`RANDOM}};
  lineBuffer_439_value = _RAND_888[7:0];
  _RAND_889 = {1{`RANDOM}};
  lineBuffer_440_grad_dir = _RAND_889[1:0];
  _RAND_890 = {1{`RANDOM}};
  lineBuffer_440_value = _RAND_890[7:0];
  _RAND_891 = {1{`RANDOM}};
  lineBuffer_441_grad_dir = _RAND_891[1:0];
  _RAND_892 = {1{`RANDOM}};
  lineBuffer_441_value = _RAND_892[7:0];
  _RAND_893 = {1{`RANDOM}};
  lineBuffer_442_grad_dir = _RAND_893[1:0];
  _RAND_894 = {1{`RANDOM}};
  lineBuffer_442_value = _RAND_894[7:0];
  _RAND_895 = {1{`RANDOM}};
  lineBuffer_443_grad_dir = _RAND_895[1:0];
  _RAND_896 = {1{`RANDOM}};
  lineBuffer_443_value = _RAND_896[7:0];
  _RAND_897 = {1{`RANDOM}};
  lineBuffer_444_grad_dir = _RAND_897[1:0];
  _RAND_898 = {1{`RANDOM}};
  lineBuffer_444_value = _RAND_898[7:0];
  _RAND_899 = {1{`RANDOM}};
  lineBuffer_445_grad_dir = _RAND_899[1:0];
  _RAND_900 = {1{`RANDOM}};
  lineBuffer_445_value = _RAND_900[7:0];
  _RAND_901 = {1{`RANDOM}};
  lineBuffer_446_grad_dir = _RAND_901[1:0];
  _RAND_902 = {1{`RANDOM}};
  lineBuffer_446_value = _RAND_902[7:0];
  _RAND_903 = {1{`RANDOM}};
  lineBuffer_447_grad_dir = _RAND_903[1:0];
  _RAND_904 = {1{`RANDOM}};
  lineBuffer_447_value = _RAND_904[7:0];
  _RAND_905 = {1{`RANDOM}};
  lineBuffer_448_grad_dir = _RAND_905[1:0];
  _RAND_906 = {1{`RANDOM}};
  lineBuffer_448_value = _RAND_906[7:0];
  _RAND_907 = {1{`RANDOM}};
  lineBuffer_449_grad_dir = _RAND_907[1:0];
  _RAND_908 = {1{`RANDOM}};
  lineBuffer_449_value = _RAND_908[7:0];
  _RAND_909 = {1{`RANDOM}};
  lineBuffer_450_grad_dir = _RAND_909[1:0];
  _RAND_910 = {1{`RANDOM}};
  lineBuffer_450_value = _RAND_910[7:0];
  _RAND_911 = {1{`RANDOM}};
  lineBuffer_451_grad_dir = _RAND_911[1:0];
  _RAND_912 = {1{`RANDOM}};
  lineBuffer_451_value = _RAND_912[7:0];
  _RAND_913 = {1{`RANDOM}};
  lineBuffer_452_grad_dir = _RAND_913[1:0];
  _RAND_914 = {1{`RANDOM}};
  lineBuffer_452_value = _RAND_914[7:0];
  _RAND_915 = {1{`RANDOM}};
  lineBuffer_453_grad_dir = _RAND_915[1:0];
  _RAND_916 = {1{`RANDOM}};
  lineBuffer_453_value = _RAND_916[7:0];
  _RAND_917 = {1{`RANDOM}};
  lineBuffer_454_grad_dir = _RAND_917[1:0];
  _RAND_918 = {1{`RANDOM}};
  lineBuffer_454_value = _RAND_918[7:0];
  _RAND_919 = {1{`RANDOM}};
  lineBuffer_455_grad_dir = _RAND_919[1:0];
  _RAND_920 = {1{`RANDOM}};
  lineBuffer_455_value = _RAND_920[7:0];
  _RAND_921 = {1{`RANDOM}};
  lineBuffer_456_grad_dir = _RAND_921[1:0];
  _RAND_922 = {1{`RANDOM}};
  lineBuffer_456_value = _RAND_922[7:0];
  _RAND_923 = {1{`RANDOM}};
  lineBuffer_457_grad_dir = _RAND_923[1:0];
  _RAND_924 = {1{`RANDOM}};
  lineBuffer_457_value = _RAND_924[7:0];
  _RAND_925 = {1{`RANDOM}};
  lineBuffer_458_grad_dir = _RAND_925[1:0];
  _RAND_926 = {1{`RANDOM}};
  lineBuffer_458_value = _RAND_926[7:0];
  _RAND_927 = {1{`RANDOM}};
  lineBuffer_459_grad_dir = _RAND_927[1:0];
  _RAND_928 = {1{`RANDOM}};
  lineBuffer_459_value = _RAND_928[7:0];
  _RAND_929 = {1{`RANDOM}};
  lineBuffer_460_grad_dir = _RAND_929[1:0];
  _RAND_930 = {1{`RANDOM}};
  lineBuffer_460_value = _RAND_930[7:0];
  _RAND_931 = {1{`RANDOM}};
  lineBuffer_461_grad_dir = _RAND_931[1:0];
  _RAND_932 = {1{`RANDOM}};
  lineBuffer_461_value = _RAND_932[7:0];
  _RAND_933 = {1{`RANDOM}};
  lineBuffer_462_grad_dir = _RAND_933[1:0];
  _RAND_934 = {1{`RANDOM}};
  lineBuffer_462_value = _RAND_934[7:0];
  _RAND_935 = {1{`RANDOM}};
  lineBuffer_463_grad_dir = _RAND_935[1:0];
  _RAND_936 = {1{`RANDOM}};
  lineBuffer_463_value = _RAND_936[7:0];
  _RAND_937 = {1{`RANDOM}};
  lineBuffer_464_grad_dir = _RAND_937[1:0];
  _RAND_938 = {1{`RANDOM}};
  lineBuffer_464_value = _RAND_938[7:0];
  _RAND_939 = {1{`RANDOM}};
  lineBuffer_465_grad_dir = _RAND_939[1:0];
  _RAND_940 = {1{`RANDOM}};
  lineBuffer_465_value = _RAND_940[7:0];
  _RAND_941 = {1{`RANDOM}};
  lineBuffer_466_grad_dir = _RAND_941[1:0];
  _RAND_942 = {1{`RANDOM}};
  lineBuffer_466_value = _RAND_942[7:0];
  _RAND_943 = {1{`RANDOM}};
  lineBuffer_467_grad_dir = _RAND_943[1:0];
  _RAND_944 = {1{`RANDOM}};
  lineBuffer_467_value = _RAND_944[7:0];
  _RAND_945 = {1{`RANDOM}};
  lineBuffer_468_grad_dir = _RAND_945[1:0];
  _RAND_946 = {1{`RANDOM}};
  lineBuffer_468_value = _RAND_946[7:0];
  _RAND_947 = {1{`RANDOM}};
  lineBuffer_469_grad_dir = _RAND_947[1:0];
  _RAND_948 = {1{`RANDOM}};
  lineBuffer_469_value = _RAND_948[7:0];
  _RAND_949 = {1{`RANDOM}};
  lineBuffer_470_grad_dir = _RAND_949[1:0];
  _RAND_950 = {1{`RANDOM}};
  lineBuffer_470_value = _RAND_950[7:0];
  _RAND_951 = {1{`RANDOM}};
  lineBuffer_471_grad_dir = _RAND_951[1:0];
  _RAND_952 = {1{`RANDOM}};
  lineBuffer_471_value = _RAND_952[7:0];
  _RAND_953 = {1{`RANDOM}};
  lineBuffer_472_grad_dir = _RAND_953[1:0];
  _RAND_954 = {1{`RANDOM}};
  lineBuffer_472_value = _RAND_954[7:0];
  _RAND_955 = {1{`RANDOM}};
  lineBuffer_473_grad_dir = _RAND_955[1:0];
  _RAND_956 = {1{`RANDOM}};
  lineBuffer_473_value = _RAND_956[7:0];
  _RAND_957 = {1{`RANDOM}};
  lineBuffer_474_grad_dir = _RAND_957[1:0];
  _RAND_958 = {1{`RANDOM}};
  lineBuffer_474_value = _RAND_958[7:0];
  _RAND_959 = {1{`RANDOM}};
  lineBuffer_475_grad_dir = _RAND_959[1:0];
  _RAND_960 = {1{`RANDOM}};
  lineBuffer_475_value = _RAND_960[7:0];
  _RAND_961 = {1{`RANDOM}};
  lineBuffer_476_grad_dir = _RAND_961[1:0];
  _RAND_962 = {1{`RANDOM}};
  lineBuffer_476_value = _RAND_962[7:0];
  _RAND_963 = {1{`RANDOM}};
  lineBuffer_477_grad_dir = _RAND_963[1:0];
  _RAND_964 = {1{`RANDOM}};
  lineBuffer_477_value = _RAND_964[7:0];
  _RAND_965 = {1{`RANDOM}};
  lineBuffer_478_grad_dir = _RAND_965[1:0];
  _RAND_966 = {1{`RANDOM}};
  lineBuffer_478_value = _RAND_966[7:0];
  _RAND_967 = {1{`RANDOM}};
  lineBuffer_479_grad_dir = _RAND_967[1:0];
  _RAND_968 = {1{`RANDOM}};
  lineBuffer_479_value = _RAND_968[7:0];
  _RAND_969 = {1{`RANDOM}};
  lineBuffer_480_grad_dir = _RAND_969[1:0];
  _RAND_970 = {1{`RANDOM}};
  lineBuffer_480_value = _RAND_970[7:0];
  _RAND_971 = {1{`RANDOM}};
  lineBuffer_481_grad_dir = _RAND_971[1:0];
  _RAND_972 = {1{`RANDOM}};
  lineBuffer_481_value = _RAND_972[7:0];
  _RAND_973 = {1{`RANDOM}};
  lineBuffer_482_grad_dir = _RAND_973[1:0];
  _RAND_974 = {1{`RANDOM}};
  lineBuffer_482_value = _RAND_974[7:0];
  _RAND_975 = {1{`RANDOM}};
  lineBuffer_483_grad_dir = _RAND_975[1:0];
  _RAND_976 = {1{`RANDOM}};
  lineBuffer_483_value = _RAND_976[7:0];
  _RAND_977 = {1{`RANDOM}};
  lineBuffer_484_grad_dir = _RAND_977[1:0];
  _RAND_978 = {1{`RANDOM}};
  lineBuffer_484_value = _RAND_978[7:0];
  _RAND_979 = {1{`RANDOM}};
  lineBuffer_485_grad_dir = _RAND_979[1:0];
  _RAND_980 = {1{`RANDOM}};
  lineBuffer_485_value = _RAND_980[7:0];
  _RAND_981 = {1{`RANDOM}};
  lineBuffer_486_grad_dir = _RAND_981[1:0];
  _RAND_982 = {1{`RANDOM}};
  lineBuffer_486_value = _RAND_982[7:0];
  _RAND_983 = {1{`RANDOM}};
  lineBuffer_487_grad_dir = _RAND_983[1:0];
  _RAND_984 = {1{`RANDOM}};
  lineBuffer_487_value = _RAND_984[7:0];
  _RAND_985 = {1{`RANDOM}};
  lineBuffer_488_grad_dir = _RAND_985[1:0];
  _RAND_986 = {1{`RANDOM}};
  lineBuffer_488_value = _RAND_986[7:0];
  _RAND_987 = {1{`RANDOM}};
  lineBuffer_489_grad_dir = _RAND_987[1:0];
  _RAND_988 = {1{`RANDOM}};
  lineBuffer_489_value = _RAND_988[7:0];
  _RAND_989 = {1{`RANDOM}};
  lineBuffer_490_grad_dir = _RAND_989[1:0];
  _RAND_990 = {1{`RANDOM}};
  lineBuffer_490_value = _RAND_990[7:0];
  _RAND_991 = {1{`RANDOM}};
  lineBuffer_491_grad_dir = _RAND_991[1:0];
  _RAND_992 = {1{`RANDOM}};
  lineBuffer_491_value = _RAND_992[7:0];
  _RAND_993 = {1{`RANDOM}};
  lineBuffer_492_grad_dir = _RAND_993[1:0];
  _RAND_994 = {1{`RANDOM}};
  lineBuffer_492_value = _RAND_994[7:0];
  _RAND_995 = {1{`RANDOM}};
  lineBuffer_493_grad_dir = _RAND_995[1:0];
  _RAND_996 = {1{`RANDOM}};
  lineBuffer_493_value = _RAND_996[7:0];
  _RAND_997 = {1{`RANDOM}};
  lineBuffer_494_grad_dir = _RAND_997[1:0];
  _RAND_998 = {1{`RANDOM}};
  lineBuffer_494_value = _RAND_998[7:0];
  _RAND_999 = {1{`RANDOM}};
  lineBuffer_495_grad_dir = _RAND_999[1:0];
  _RAND_1000 = {1{`RANDOM}};
  lineBuffer_495_value = _RAND_1000[7:0];
  _RAND_1001 = {1{`RANDOM}};
  lineBuffer_496_grad_dir = _RAND_1001[1:0];
  _RAND_1002 = {1{`RANDOM}};
  lineBuffer_496_value = _RAND_1002[7:0];
  _RAND_1003 = {1{`RANDOM}};
  lineBuffer_497_grad_dir = _RAND_1003[1:0];
  _RAND_1004 = {1{`RANDOM}};
  lineBuffer_497_value = _RAND_1004[7:0];
  _RAND_1005 = {1{`RANDOM}};
  lineBuffer_498_grad_dir = _RAND_1005[1:0];
  _RAND_1006 = {1{`RANDOM}};
  lineBuffer_498_value = _RAND_1006[7:0];
  _RAND_1007 = {1{`RANDOM}};
  lineBuffer_499_grad_dir = _RAND_1007[1:0];
  _RAND_1008 = {1{`RANDOM}};
  lineBuffer_499_value = _RAND_1008[7:0];
  _RAND_1009 = {1{`RANDOM}};
  lineBuffer_500_grad_dir = _RAND_1009[1:0];
  _RAND_1010 = {1{`RANDOM}};
  lineBuffer_500_value = _RAND_1010[7:0];
  _RAND_1011 = {1{`RANDOM}};
  lineBuffer_501_grad_dir = _RAND_1011[1:0];
  _RAND_1012 = {1{`RANDOM}};
  lineBuffer_501_value = _RAND_1012[7:0];
  _RAND_1013 = {1{`RANDOM}};
  lineBuffer_502_grad_dir = _RAND_1013[1:0];
  _RAND_1014 = {1{`RANDOM}};
  lineBuffer_502_value = _RAND_1014[7:0];
  _RAND_1015 = {1{`RANDOM}};
  lineBuffer_503_grad_dir = _RAND_1015[1:0];
  _RAND_1016 = {1{`RANDOM}};
  lineBuffer_503_value = _RAND_1016[7:0];
  _RAND_1017 = {1{`RANDOM}};
  lineBuffer_504_grad_dir = _RAND_1017[1:0];
  _RAND_1018 = {1{`RANDOM}};
  lineBuffer_504_value = _RAND_1018[7:0];
  _RAND_1019 = {1{`RANDOM}};
  lineBuffer_505_grad_dir = _RAND_1019[1:0];
  _RAND_1020 = {1{`RANDOM}};
  lineBuffer_505_value = _RAND_1020[7:0];
  _RAND_1021 = {1{`RANDOM}};
  lineBuffer_506_grad_dir = _RAND_1021[1:0];
  _RAND_1022 = {1{`RANDOM}};
  lineBuffer_506_value = _RAND_1022[7:0];
  _RAND_1023 = {1{`RANDOM}};
  lineBuffer_507_grad_dir = _RAND_1023[1:0];
  _RAND_1024 = {1{`RANDOM}};
  lineBuffer_507_value = _RAND_1024[7:0];
  _RAND_1025 = {1{`RANDOM}};
  lineBuffer_508_grad_dir = _RAND_1025[1:0];
  _RAND_1026 = {1{`RANDOM}};
  lineBuffer_508_value = _RAND_1026[7:0];
  _RAND_1027 = {1{`RANDOM}};
  lineBuffer_509_grad_dir = _RAND_1027[1:0];
  _RAND_1028 = {1{`RANDOM}};
  lineBuffer_509_value = _RAND_1028[7:0];
  _RAND_1029 = {1{`RANDOM}};
  lineBuffer_510_grad_dir = _RAND_1029[1:0];
  _RAND_1030 = {1{`RANDOM}};
  lineBuffer_510_value = _RAND_1030[7:0];
  _RAND_1031 = {1{`RANDOM}};
  lineBuffer_511_grad_dir = _RAND_1031[1:0];
  _RAND_1032 = {1{`RANDOM}};
  lineBuffer_511_value = _RAND_1032[7:0];
  _RAND_1033 = {1{`RANDOM}};
  lineBuffer_512_value = _RAND_1033[7:0];
  _RAND_1034 = {1{`RANDOM}};
  lineBuffer_513_value = _RAND_1034[7:0];
  _RAND_1035 = {1{`RANDOM}};
  lineBuffer_514_value = _RAND_1035[7:0];
  _RAND_1036 = {1{`RANDOM}};
  lineBuffer_515_value = _RAND_1036[7:0];
  _RAND_1037 = {1{`RANDOM}};
  lineBuffer_516_value = _RAND_1037[7:0];
  _RAND_1038 = {1{`RANDOM}};
  lineBuffer_517_value = _RAND_1038[7:0];
  _RAND_1039 = {1{`RANDOM}};
  lineBuffer_518_value = _RAND_1039[7:0];
  _RAND_1040 = {1{`RANDOM}};
  lineBuffer_519_value = _RAND_1040[7:0];
  _RAND_1041 = {1{`RANDOM}};
  lineBuffer_520_value = _RAND_1041[7:0];
  _RAND_1042 = {1{`RANDOM}};
  lineBuffer_521_value = _RAND_1042[7:0];
  _RAND_1043 = {1{`RANDOM}};
  lineBuffer_522_value = _RAND_1043[7:0];
  _RAND_1044 = {1{`RANDOM}};
  lineBuffer_523_value = _RAND_1044[7:0];
  _RAND_1045 = {1{`RANDOM}};
  lineBuffer_524_value = _RAND_1045[7:0];
  _RAND_1046 = {1{`RANDOM}};
  lineBuffer_525_value = _RAND_1046[7:0];
  _RAND_1047 = {1{`RANDOM}};
  lineBuffer_526_value = _RAND_1047[7:0];
  _RAND_1048 = {1{`RANDOM}};
  lineBuffer_527_value = _RAND_1048[7:0];
  _RAND_1049 = {1{`RANDOM}};
  lineBuffer_528_value = _RAND_1049[7:0];
  _RAND_1050 = {1{`RANDOM}};
  lineBuffer_529_value = _RAND_1050[7:0];
  _RAND_1051 = {1{`RANDOM}};
  lineBuffer_530_value = _RAND_1051[7:0];
  _RAND_1052 = {1{`RANDOM}};
  lineBuffer_531_value = _RAND_1052[7:0];
  _RAND_1053 = {1{`RANDOM}};
  lineBuffer_532_value = _RAND_1053[7:0];
  _RAND_1054 = {1{`RANDOM}};
  lineBuffer_533_value = _RAND_1054[7:0];
  _RAND_1055 = {1{`RANDOM}};
  lineBuffer_534_value = _RAND_1055[7:0];
  _RAND_1056 = {1{`RANDOM}};
  lineBuffer_535_value = _RAND_1056[7:0];
  _RAND_1057 = {1{`RANDOM}};
  lineBuffer_536_value = _RAND_1057[7:0];
  _RAND_1058 = {1{`RANDOM}};
  lineBuffer_537_value = _RAND_1058[7:0];
  _RAND_1059 = {1{`RANDOM}};
  lineBuffer_538_value = _RAND_1059[7:0];
  _RAND_1060 = {1{`RANDOM}};
  lineBuffer_539_value = _RAND_1060[7:0];
  _RAND_1061 = {1{`RANDOM}};
  lineBuffer_540_value = _RAND_1061[7:0];
  _RAND_1062 = {1{`RANDOM}};
  lineBuffer_541_value = _RAND_1062[7:0];
  _RAND_1063 = {1{`RANDOM}};
  lineBuffer_542_value = _RAND_1063[7:0];
  _RAND_1064 = {1{`RANDOM}};
  lineBuffer_543_value = _RAND_1064[7:0];
  _RAND_1065 = {1{`RANDOM}};
  lineBuffer_544_value = _RAND_1065[7:0];
  _RAND_1066 = {1{`RANDOM}};
  lineBuffer_545_value = _RAND_1066[7:0];
  _RAND_1067 = {1{`RANDOM}};
  lineBuffer_546_value = _RAND_1067[7:0];
  _RAND_1068 = {1{`RANDOM}};
  lineBuffer_547_value = _RAND_1068[7:0];
  _RAND_1069 = {1{`RANDOM}};
  lineBuffer_548_value = _RAND_1069[7:0];
  _RAND_1070 = {1{`RANDOM}};
  lineBuffer_549_value = _RAND_1070[7:0];
  _RAND_1071 = {1{`RANDOM}};
  lineBuffer_550_value = _RAND_1071[7:0];
  _RAND_1072 = {1{`RANDOM}};
  lineBuffer_551_value = _RAND_1072[7:0];
  _RAND_1073 = {1{`RANDOM}};
  lineBuffer_552_value = _RAND_1073[7:0];
  _RAND_1074 = {1{`RANDOM}};
  lineBuffer_553_value = _RAND_1074[7:0];
  _RAND_1075 = {1{`RANDOM}};
  lineBuffer_554_value = _RAND_1075[7:0];
  _RAND_1076 = {1{`RANDOM}};
  lineBuffer_555_value = _RAND_1076[7:0];
  _RAND_1077 = {1{`RANDOM}};
  lineBuffer_556_value = _RAND_1077[7:0];
  _RAND_1078 = {1{`RANDOM}};
  lineBuffer_557_value = _RAND_1078[7:0];
  _RAND_1079 = {1{`RANDOM}};
  lineBuffer_558_value = _RAND_1079[7:0];
  _RAND_1080 = {1{`RANDOM}};
  lineBuffer_559_value = _RAND_1080[7:0];
  _RAND_1081 = {1{`RANDOM}};
  lineBuffer_560_value = _RAND_1081[7:0];
  _RAND_1082 = {1{`RANDOM}};
  lineBuffer_561_value = _RAND_1082[7:0];
  _RAND_1083 = {1{`RANDOM}};
  lineBuffer_562_value = _RAND_1083[7:0];
  _RAND_1084 = {1{`RANDOM}};
  lineBuffer_563_value = _RAND_1084[7:0];
  _RAND_1085 = {1{`RANDOM}};
  lineBuffer_564_value = _RAND_1085[7:0];
  _RAND_1086 = {1{`RANDOM}};
  lineBuffer_565_value = _RAND_1086[7:0];
  _RAND_1087 = {1{`RANDOM}};
  lineBuffer_566_value = _RAND_1087[7:0];
  _RAND_1088 = {1{`RANDOM}};
  lineBuffer_567_value = _RAND_1088[7:0];
  _RAND_1089 = {1{`RANDOM}};
  lineBuffer_568_value = _RAND_1089[7:0];
  _RAND_1090 = {1{`RANDOM}};
  lineBuffer_569_value = _RAND_1090[7:0];
  _RAND_1091 = {1{`RANDOM}};
  lineBuffer_570_value = _RAND_1091[7:0];
  _RAND_1092 = {1{`RANDOM}};
  lineBuffer_571_value = _RAND_1092[7:0];
  _RAND_1093 = {1{`RANDOM}};
  lineBuffer_572_value = _RAND_1093[7:0];
  _RAND_1094 = {1{`RANDOM}};
  lineBuffer_573_value = _RAND_1094[7:0];
  _RAND_1095 = {1{`RANDOM}};
  lineBuffer_574_value = _RAND_1095[7:0];
  _RAND_1096 = {1{`RANDOM}};
  lineBuffer_575_value = _RAND_1096[7:0];
  _RAND_1097 = {1{`RANDOM}};
  lineBuffer_576_value = _RAND_1097[7:0];
  _RAND_1098 = {1{`RANDOM}};
  lineBuffer_577_value = _RAND_1098[7:0];
  _RAND_1099 = {1{`RANDOM}};
  lineBuffer_578_value = _RAND_1099[7:0];
  _RAND_1100 = {1{`RANDOM}};
  lineBuffer_579_value = _RAND_1100[7:0];
  _RAND_1101 = {1{`RANDOM}};
  lineBuffer_580_value = _RAND_1101[7:0];
  _RAND_1102 = {1{`RANDOM}};
  lineBuffer_581_value = _RAND_1102[7:0];
  _RAND_1103 = {1{`RANDOM}};
  lineBuffer_582_value = _RAND_1103[7:0];
  _RAND_1104 = {1{`RANDOM}};
  lineBuffer_583_value = _RAND_1104[7:0];
  _RAND_1105 = {1{`RANDOM}};
  lineBuffer_584_value = _RAND_1105[7:0];
  _RAND_1106 = {1{`RANDOM}};
  lineBuffer_585_value = _RAND_1106[7:0];
  _RAND_1107 = {1{`RANDOM}};
  lineBuffer_586_value = _RAND_1107[7:0];
  _RAND_1108 = {1{`RANDOM}};
  lineBuffer_587_value = _RAND_1108[7:0];
  _RAND_1109 = {1{`RANDOM}};
  lineBuffer_588_value = _RAND_1109[7:0];
  _RAND_1110 = {1{`RANDOM}};
  lineBuffer_589_value = _RAND_1110[7:0];
  _RAND_1111 = {1{`RANDOM}};
  lineBuffer_590_value = _RAND_1111[7:0];
  _RAND_1112 = {1{`RANDOM}};
  lineBuffer_591_value = _RAND_1112[7:0];
  _RAND_1113 = {1{`RANDOM}};
  lineBuffer_592_value = _RAND_1113[7:0];
  _RAND_1114 = {1{`RANDOM}};
  lineBuffer_593_value = _RAND_1114[7:0];
  _RAND_1115 = {1{`RANDOM}};
  lineBuffer_594_value = _RAND_1115[7:0];
  _RAND_1116 = {1{`RANDOM}};
  lineBuffer_595_value = _RAND_1116[7:0];
  _RAND_1117 = {1{`RANDOM}};
  lineBuffer_596_value = _RAND_1117[7:0];
  _RAND_1118 = {1{`RANDOM}};
  lineBuffer_597_value = _RAND_1118[7:0];
  _RAND_1119 = {1{`RANDOM}};
  lineBuffer_598_value = _RAND_1119[7:0];
  _RAND_1120 = {1{`RANDOM}};
  lineBuffer_599_value = _RAND_1120[7:0];
  _RAND_1121 = {1{`RANDOM}};
  lineBuffer_600_value = _RAND_1121[7:0];
  _RAND_1122 = {1{`RANDOM}};
  lineBuffer_601_value = _RAND_1122[7:0];
  _RAND_1123 = {1{`RANDOM}};
  lineBuffer_602_value = _RAND_1123[7:0];
  _RAND_1124 = {1{`RANDOM}};
  lineBuffer_603_value = _RAND_1124[7:0];
  _RAND_1125 = {1{`RANDOM}};
  lineBuffer_604_value = _RAND_1125[7:0];
  _RAND_1126 = {1{`RANDOM}};
  lineBuffer_605_value = _RAND_1126[7:0];
  _RAND_1127 = {1{`RANDOM}};
  lineBuffer_606_value = _RAND_1127[7:0];
  _RAND_1128 = {1{`RANDOM}};
  lineBuffer_607_value = _RAND_1128[7:0];
  _RAND_1129 = {1{`RANDOM}};
  lineBuffer_608_value = _RAND_1129[7:0];
  _RAND_1130 = {1{`RANDOM}};
  lineBuffer_609_value = _RAND_1130[7:0];
  _RAND_1131 = {1{`RANDOM}};
  lineBuffer_610_value = _RAND_1131[7:0];
  _RAND_1132 = {1{`RANDOM}};
  lineBuffer_611_value = _RAND_1132[7:0];
  _RAND_1133 = {1{`RANDOM}};
  lineBuffer_612_value = _RAND_1133[7:0];
  _RAND_1134 = {1{`RANDOM}};
  lineBuffer_613_value = _RAND_1134[7:0];
  _RAND_1135 = {1{`RANDOM}};
  lineBuffer_614_value = _RAND_1135[7:0];
  _RAND_1136 = {1{`RANDOM}};
  lineBuffer_615_value = _RAND_1136[7:0];
  _RAND_1137 = {1{`RANDOM}};
  lineBuffer_616_value = _RAND_1137[7:0];
  _RAND_1138 = {1{`RANDOM}};
  lineBuffer_617_value = _RAND_1138[7:0];
  _RAND_1139 = {1{`RANDOM}};
  lineBuffer_618_value = _RAND_1139[7:0];
  _RAND_1140 = {1{`RANDOM}};
  lineBuffer_619_value = _RAND_1140[7:0];
  _RAND_1141 = {1{`RANDOM}};
  lineBuffer_620_value = _RAND_1141[7:0];
  _RAND_1142 = {1{`RANDOM}};
  lineBuffer_621_value = _RAND_1142[7:0];
  _RAND_1143 = {1{`RANDOM}};
  lineBuffer_622_value = _RAND_1143[7:0];
  _RAND_1144 = {1{`RANDOM}};
  lineBuffer_623_value = _RAND_1144[7:0];
  _RAND_1145 = {1{`RANDOM}};
  lineBuffer_624_value = _RAND_1145[7:0];
  _RAND_1146 = {1{`RANDOM}};
  lineBuffer_625_value = _RAND_1146[7:0];
  _RAND_1147 = {1{`RANDOM}};
  lineBuffer_626_value = _RAND_1147[7:0];
  _RAND_1148 = {1{`RANDOM}};
  lineBuffer_627_value = _RAND_1148[7:0];
  _RAND_1149 = {1{`RANDOM}};
  lineBuffer_628_value = _RAND_1149[7:0];
  _RAND_1150 = {1{`RANDOM}};
  lineBuffer_629_value = _RAND_1150[7:0];
  _RAND_1151 = {1{`RANDOM}};
  lineBuffer_630_value = _RAND_1151[7:0];
  _RAND_1152 = {1{`RANDOM}};
  lineBuffer_631_value = _RAND_1152[7:0];
  _RAND_1153 = {1{`RANDOM}};
  lineBuffer_632_value = _RAND_1153[7:0];
  _RAND_1154 = {1{`RANDOM}};
  lineBuffer_633_value = _RAND_1154[7:0];
  _RAND_1155 = {1{`RANDOM}};
  lineBuffer_634_value = _RAND_1155[7:0];
  _RAND_1156 = {1{`RANDOM}};
  lineBuffer_635_value = _RAND_1156[7:0];
  _RAND_1157 = {1{`RANDOM}};
  lineBuffer_636_value = _RAND_1157[7:0];
  _RAND_1158 = {1{`RANDOM}};
  lineBuffer_637_value = _RAND_1158[7:0];
  _RAND_1159 = {1{`RANDOM}};
  lineBuffer_638_value = _RAND_1159[7:0];
  _RAND_1160 = {1{`RANDOM}};
  lineBuffer_639_value = _RAND_1160[7:0];
  _RAND_1161 = {1{`RANDOM}};
  lineBuffer_640_value = _RAND_1161[7:0];
  _RAND_1162 = {1{`RANDOM}};
  lineBuffer_641_value = _RAND_1162[7:0];
  _RAND_1163 = {1{`RANDOM}};
  lineBuffer_642_value = _RAND_1163[7:0];
  _RAND_1164 = {1{`RANDOM}};
  lineBuffer_643_value = _RAND_1164[7:0];
  _RAND_1165 = {1{`RANDOM}};
  lineBuffer_644_value = _RAND_1165[7:0];
  _RAND_1166 = {1{`RANDOM}};
  lineBuffer_645_value = _RAND_1166[7:0];
  _RAND_1167 = {1{`RANDOM}};
  lineBuffer_646_value = _RAND_1167[7:0];
  _RAND_1168 = {1{`RANDOM}};
  lineBuffer_647_value = _RAND_1168[7:0];
  _RAND_1169 = {1{`RANDOM}};
  lineBuffer_648_value = _RAND_1169[7:0];
  _RAND_1170 = {1{`RANDOM}};
  lineBuffer_649_value = _RAND_1170[7:0];
  _RAND_1171 = {1{`RANDOM}};
  lineBuffer_650_value = _RAND_1171[7:0];
  _RAND_1172 = {1{`RANDOM}};
  lineBuffer_651_value = _RAND_1172[7:0];
  _RAND_1173 = {1{`RANDOM}};
  lineBuffer_652_value = _RAND_1173[7:0];
  _RAND_1174 = {1{`RANDOM}};
  lineBuffer_653_value = _RAND_1174[7:0];
  _RAND_1175 = {1{`RANDOM}};
  lineBuffer_654_value = _RAND_1175[7:0];
  _RAND_1176 = {1{`RANDOM}};
  lineBuffer_655_value = _RAND_1176[7:0];
  _RAND_1177 = {1{`RANDOM}};
  lineBuffer_656_value = _RAND_1177[7:0];
  _RAND_1178 = {1{`RANDOM}};
  lineBuffer_657_value = _RAND_1178[7:0];
  _RAND_1179 = {1{`RANDOM}};
  lineBuffer_658_value = _RAND_1179[7:0];
  _RAND_1180 = {1{`RANDOM}};
  lineBuffer_659_value = _RAND_1180[7:0];
  _RAND_1181 = {1{`RANDOM}};
  lineBuffer_660_value = _RAND_1181[7:0];
  _RAND_1182 = {1{`RANDOM}};
  lineBuffer_661_value = _RAND_1182[7:0];
  _RAND_1183 = {1{`RANDOM}};
  lineBuffer_662_value = _RAND_1183[7:0];
  _RAND_1184 = {1{`RANDOM}};
  lineBuffer_663_value = _RAND_1184[7:0];
  _RAND_1185 = {1{`RANDOM}};
  lineBuffer_664_value = _RAND_1185[7:0];
  _RAND_1186 = {1{`RANDOM}};
  lineBuffer_665_value = _RAND_1186[7:0];
  _RAND_1187 = {1{`RANDOM}};
  lineBuffer_666_value = _RAND_1187[7:0];
  _RAND_1188 = {1{`RANDOM}};
  lineBuffer_667_value = _RAND_1188[7:0];
  _RAND_1189 = {1{`RANDOM}};
  lineBuffer_668_value = _RAND_1189[7:0];
  _RAND_1190 = {1{`RANDOM}};
  lineBuffer_669_value = _RAND_1190[7:0];
  _RAND_1191 = {1{`RANDOM}};
  lineBuffer_670_value = _RAND_1191[7:0];
  _RAND_1192 = {1{`RANDOM}};
  lineBuffer_671_value = _RAND_1192[7:0];
  _RAND_1193 = {1{`RANDOM}};
  lineBuffer_672_value = _RAND_1193[7:0];
  _RAND_1194 = {1{`RANDOM}};
  lineBuffer_673_value = _RAND_1194[7:0];
  _RAND_1195 = {1{`RANDOM}};
  lineBuffer_674_value = _RAND_1195[7:0];
  _RAND_1196 = {1{`RANDOM}};
  lineBuffer_675_value = _RAND_1196[7:0];
  _RAND_1197 = {1{`RANDOM}};
  lineBuffer_676_value = _RAND_1197[7:0];
  _RAND_1198 = {1{`RANDOM}};
  lineBuffer_677_value = _RAND_1198[7:0];
  _RAND_1199 = {1{`RANDOM}};
  lineBuffer_678_value = _RAND_1199[7:0];
  _RAND_1200 = {1{`RANDOM}};
  lineBuffer_679_value = _RAND_1200[7:0];
  _RAND_1201 = {1{`RANDOM}};
  lineBuffer_680_value = _RAND_1201[7:0];
  _RAND_1202 = {1{`RANDOM}};
  lineBuffer_681_value = _RAND_1202[7:0];
  _RAND_1203 = {1{`RANDOM}};
  lineBuffer_682_value = _RAND_1203[7:0];
  _RAND_1204 = {1{`RANDOM}};
  lineBuffer_683_value = _RAND_1204[7:0];
  _RAND_1205 = {1{`RANDOM}};
  lineBuffer_684_value = _RAND_1205[7:0];
  _RAND_1206 = {1{`RANDOM}};
  lineBuffer_685_value = _RAND_1206[7:0];
  _RAND_1207 = {1{`RANDOM}};
  lineBuffer_686_value = _RAND_1207[7:0];
  _RAND_1208 = {1{`RANDOM}};
  lineBuffer_687_value = _RAND_1208[7:0];
  _RAND_1209 = {1{`RANDOM}};
  lineBuffer_688_value = _RAND_1209[7:0];
  _RAND_1210 = {1{`RANDOM}};
  lineBuffer_689_value = _RAND_1210[7:0];
  _RAND_1211 = {1{`RANDOM}};
  lineBuffer_690_value = _RAND_1211[7:0];
  _RAND_1212 = {1{`RANDOM}};
  lineBuffer_691_value = _RAND_1212[7:0];
  _RAND_1213 = {1{`RANDOM}};
  lineBuffer_692_value = _RAND_1213[7:0];
  _RAND_1214 = {1{`RANDOM}};
  lineBuffer_693_value = _RAND_1214[7:0];
  _RAND_1215 = {1{`RANDOM}};
  lineBuffer_694_value = _RAND_1215[7:0];
  _RAND_1216 = {1{`RANDOM}};
  lineBuffer_695_value = _RAND_1216[7:0];
  _RAND_1217 = {1{`RANDOM}};
  lineBuffer_696_value = _RAND_1217[7:0];
  _RAND_1218 = {1{`RANDOM}};
  lineBuffer_697_value = _RAND_1218[7:0];
  _RAND_1219 = {1{`RANDOM}};
  lineBuffer_698_value = _RAND_1219[7:0];
  _RAND_1220 = {1{`RANDOM}};
  lineBuffer_699_value = _RAND_1220[7:0];
  _RAND_1221 = {1{`RANDOM}};
  lineBuffer_700_value = _RAND_1221[7:0];
  _RAND_1222 = {1{`RANDOM}};
  lineBuffer_701_value = _RAND_1222[7:0];
  _RAND_1223 = {1{`RANDOM}};
  lineBuffer_702_value = _RAND_1223[7:0];
  _RAND_1224 = {1{`RANDOM}};
  lineBuffer_703_value = _RAND_1224[7:0];
  _RAND_1225 = {1{`RANDOM}};
  lineBuffer_704_value = _RAND_1225[7:0];
  _RAND_1226 = {1{`RANDOM}};
  lineBuffer_705_value = _RAND_1226[7:0];
  _RAND_1227 = {1{`RANDOM}};
  lineBuffer_706_value = _RAND_1227[7:0];
  _RAND_1228 = {1{`RANDOM}};
  lineBuffer_707_value = _RAND_1228[7:0];
  _RAND_1229 = {1{`RANDOM}};
  lineBuffer_708_value = _RAND_1229[7:0];
  _RAND_1230 = {1{`RANDOM}};
  lineBuffer_709_value = _RAND_1230[7:0];
  _RAND_1231 = {1{`RANDOM}};
  lineBuffer_710_value = _RAND_1231[7:0];
  _RAND_1232 = {1{`RANDOM}};
  lineBuffer_711_value = _RAND_1232[7:0];
  _RAND_1233 = {1{`RANDOM}};
  lineBuffer_712_value = _RAND_1233[7:0];
  _RAND_1234 = {1{`RANDOM}};
  lineBuffer_713_value = _RAND_1234[7:0];
  _RAND_1235 = {1{`RANDOM}};
  lineBuffer_714_value = _RAND_1235[7:0];
  _RAND_1236 = {1{`RANDOM}};
  lineBuffer_715_value = _RAND_1236[7:0];
  _RAND_1237 = {1{`RANDOM}};
  lineBuffer_716_value = _RAND_1237[7:0];
  _RAND_1238 = {1{`RANDOM}};
  lineBuffer_717_value = _RAND_1238[7:0];
  _RAND_1239 = {1{`RANDOM}};
  lineBuffer_718_value = _RAND_1239[7:0];
  _RAND_1240 = {1{`RANDOM}};
  lineBuffer_719_value = _RAND_1240[7:0];
  _RAND_1241 = {1{`RANDOM}};
  lineBuffer_720_value = _RAND_1241[7:0];
  _RAND_1242 = {1{`RANDOM}};
  lineBuffer_721_value = _RAND_1242[7:0];
  _RAND_1243 = {1{`RANDOM}};
  lineBuffer_722_value = _RAND_1243[7:0];
  _RAND_1244 = {1{`RANDOM}};
  lineBuffer_723_value = _RAND_1244[7:0];
  _RAND_1245 = {1{`RANDOM}};
  lineBuffer_724_value = _RAND_1245[7:0];
  _RAND_1246 = {1{`RANDOM}};
  lineBuffer_725_value = _RAND_1246[7:0];
  _RAND_1247 = {1{`RANDOM}};
  lineBuffer_726_value = _RAND_1247[7:0];
  _RAND_1248 = {1{`RANDOM}};
  lineBuffer_727_value = _RAND_1248[7:0];
  _RAND_1249 = {1{`RANDOM}};
  lineBuffer_728_value = _RAND_1249[7:0];
  _RAND_1250 = {1{`RANDOM}};
  lineBuffer_729_value = _RAND_1250[7:0];
  _RAND_1251 = {1{`RANDOM}};
  lineBuffer_730_value = _RAND_1251[7:0];
  _RAND_1252 = {1{`RANDOM}};
  lineBuffer_731_value = _RAND_1252[7:0];
  _RAND_1253 = {1{`RANDOM}};
  lineBuffer_732_value = _RAND_1253[7:0];
  _RAND_1254 = {1{`RANDOM}};
  lineBuffer_733_value = _RAND_1254[7:0];
  _RAND_1255 = {1{`RANDOM}};
  lineBuffer_734_value = _RAND_1255[7:0];
  _RAND_1256 = {1{`RANDOM}};
  lineBuffer_735_value = _RAND_1256[7:0];
  _RAND_1257 = {1{`RANDOM}};
  lineBuffer_736_value = _RAND_1257[7:0];
  _RAND_1258 = {1{`RANDOM}};
  lineBuffer_737_value = _RAND_1258[7:0];
  _RAND_1259 = {1{`RANDOM}};
  lineBuffer_738_value = _RAND_1259[7:0];
  _RAND_1260 = {1{`RANDOM}};
  lineBuffer_739_value = _RAND_1260[7:0];
  _RAND_1261 = {1{`RANDOM}};
  lineBuffer_740_value = _RAND_1261[7:0];
  _RAND_1262 = {1{`RANDOM}};
  lineBuffer_741_value = _RAND_1262[7:0];
  _RAND_1263 = {1{`RANDOM}};
  lineBuffer_742_value = _RAND_1263[7:0];
  _RAND_1264 = {1{`RANDOM}};
  lineBuffer_743_value = _RAND_1264[7:0];
  _RAND_1265 = {1{`RANDOM}};
  lineBuffer_744_value = _RAND_1265[7:0];
  _RAND_1266 = {1{`RANDOM}};
  lineBuffer_745_value = _RAND_1266[7:0];
  _RAND_1267 = {1{`RANDOM}};
  lineBuffer_746_value = _RAND_1267[7:0];
  _RAND_1268 = {1{`RANDOM}};
  lineBuffer_747_value = _RAND_1268[7:0];
  _RAND_1269 = {1{`RANDOM}};
  lineBuffer_748_value = _RAND_1269[7:0];
  _RAND_1270 = {1{`RANDOM}};
  lineBuffer_749_value = _RAND_1270[7:0];
  _RAND_1271 = {1{`RANDOM}};
  lineBuffer_750_value = _RAND_1271[7:0];
  _RAND_1272 = {1{`RANDOM}};
  lineBuffer_751_value = _RAND_1272[7:0];
  _RAND_1273 = {1{`RANDOM}};
  lineBuffer_752_value = _RAND_1273[7:0];
  _RAND_1274 = {1{`RANDOM}};
  lineBuffer_753_value = _RAND_1274[7:0];
  _RAND_1275 = {1{`RANDOM}};
  lineBuffer_754_value = _RAND_1275[7:0];
  _RAND_1276 = {1{`RANDOM}};
  lineBuffer_755_value = _RAND_1276[7:0];
  _RAND_1277 = {1{`RANDOM}};
  lineBuffer_756_value = _RAND_1277[7:0];
  _RAND_1278 = {1{`RANDOM}};
  lineBuffer_757_value = _RAND_1278[7:0];
  _RAND_1279 = {1{`RANDOM}};
  lineBuffer_758_value = _RAND_1279[7:0];
  _RAND_1280 = {1{`RANDOM}};
  lineBuffer_759_value = _RAND_1280[7:0];
  _RAND_1281 = {1{`RANDOM}};
  lineBuffer_760_value = _RAND_1281[7:0];
  _RAND_1282 = {1{`RANDOM}};
  lineBuffer_761_value = _RAND_1282[7:0];
  _RAND_1283 = {1{`RANDOM}};
  lineBuffer_762_value = _RAND_1283[7:0];
  _RAND_1284 = {1{`RANDOM}};
  lineBuffer_763_value = _RAND_1284[7:0];
  _RAND_1285 = {1{`RANDOM}};
  lineBuffer_764_value = _RAND_1285[7:0];
  _RAND_1286 = {1{`RANDOM}};
  lineBuffer_765_value = _RAND_1286[7:0];
  _RAND_1287 = {1{`RANDOM}};
  lineBuffer_766_value = _RAND_1287[7:0];
  _RAND_1288 = {1{`RANDOM}};
  lineBuffer_767_value = _RAND_1288[7:0];
  _RAND_1289 = {1{`RANDOM}};
  windowBuffer_0_value = _RAND_1289[7:0];
  _RAND_1290 = {1{`RANDOM}};
  windowBuffer_1_value = _RAND_1290[7:0];
  _RAND_1291 = {1{`RANDOM}};
  windowBuffer_2_value = _RAND_1291[7:0];
  _RAND_1292 = {1{`RANDOM}};
  windowBuffer_3_value = _RAND_1292[7:0];
  _RAND_1293 = {1{`RANDOM}};
  windowBuffer_4_grad_dir = _RAND_1293[1:0];
  _RAND_1294 = {1{`RANDOM}};
  windowBuffer_4_value = _RAND_1294[7:0];
  _RAND_1295 = {1{`RANDOM}};
  windowBuffer_5_grad_dir = _RAND_1295[1:0];
  _RAND_1296 = {1{`RANDOM}};
  windowBuffer_5_value = _RAND_1296[7:0];
  _RAND_1297 = {1{`RANDOM}};
  windowBuffer_6_value = _RAND_1297[7:0];
  _RAND_1298 = {1{`RANDOM}};
  windowBuffer_7_value = _RAND_1298[7:0];
  _RAND_1299 = {1{`RANDOM}};
  windowBuffer_8_value = _RAND_1299[7:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      stateReg <= 2'h0;
    end else if (_T) begin
      if (io_enq_valid) begin
        stateReg <= 2'h1;
      end
    end else if (_T_1) begin
      if (_T_3) begin
        stateReg <= 2'h0;
      end else if (_T_4) begin
        stateReg <= 2'h1;
      end else if (_T_6) begin
        stateReg <= 2'h2;
      end
    end else if (_T_7) begin
      if (io_deq_ready) begin
        stateReg <= 2'h1;
      end
    end else if (_T_8) begin
      stateReg <= 2'h0;
    end
    if (_T) begin
      if (io_enq_valid) begin
        dataReg_grad_dir <= io_enq_bits_grad_dir;
      end
    end else if (_T_1) begin
      if (!(_T_3)) begin
        if (_T_4) begin
          dataReg_grad_dir <= io_enq_bits_grad_dir;
        end
      end
    end else if (_T_7) begin
      if (io_deq_ready) begin
        dataReg_grad_dir <= shadowReg_grad_dir;
      end
    end
    if (_T) begin
      if (io_enq_valid) begin
        dataReg_value <= io_enq_bits_value;
      end
    end else if (_T_1) begin
      if (!(_T_3)) begin
        if (_T_4) begin
          dataReg_value <= io_enq_bits_value;
        end
      end
    end else if (_T_7) begin
      if (io_deq_ready) begin
        dataReg_value <= shadowReg_value;
      end
    end
    if (!(_T)) begin
      if (_T_1) begin
        if (!(_T_3)) begin
          if (!(_T_4)) begin
            if (_T_6) begin
              shadowReg_grad_dir <= io_enq_bits_grad_dir;
            end
          end
        end
      end
    end
    if (!(_T)) begin
      if (_T_1) begin
        if (!(_T_3)) begin
          if (!(_T_4)) begin
            if (_T_6) begin
              shadowReg_value <= io_enq_bits_value;
            end
          end
        end
      end
    end
    if (_T) begin
      userReg <= io_enq_user;
    end else if (_T_1) begin
      if (_T_3) begin
        userReg <= io_enq_user;
      end else if (_T_4) begin
        userReg <= io_enq_user;
      end
    end else if (_T_7) begin
      if (io_deq_ready) begin
        userReg <= shadowUserReg;
      end
    end
    if (!(_T)) begin
      if (_T_1) begin
        if (!(_T_3)) begin
          if (!(_T_4)) begin
            if (_T_6) begin
              shadowUserReg <= io_enq_user;
            end
          end
        end
      end
    end
    if (_T) begin
      if (io_enq_valid) begin
        lastReg <= io_enq_last;
      end
    end else if (_T_1) begin
      if (!(_T_3)) begin
        if (_T_4) begin
          lastReg <= io_enq_last;
        end
      end
    end else if (_T_7) begin
      if (io_deq_ready) begin
        lastReg <= shadowLastReg;
      end
    end
    if (!(_T)) begin
      if (_T_1) begin
        if (!(_T_3)) begin
          if (!(_T_4)) begin
            if (_T_6) begin
              shadowLastReg <= io_enq_last;
            end
          end
        end
      end
    end
    if (sel) begin
      lineBuffer_0_grad_dir <= dataReg_grad_dir;
    end
    if (sel) begin
      lineBuffer_0_value <= dataReg_value;
    end
    if (sel) begin
      lineBuffer_1_grad_dir <= lineBuffer_0_grad_dir;
    end
    if (sel) begin
      lineBuffer_1_value <= lineBuffer_0_value;
    end
    if (sel) begin
      lineBuffer_2_grad_dir <= lineBuffer_1_grad_dir;
    end
    if (sel) begin
      lineBuffer_2_value <= lineBuffer_1_value;
    end
    if (sel) begin
      lineBuffer_3_grad_dir <= lineBuffer_2_grad_dir;
    end
    if (sel) begin
      lineBuffer_3_value <= lineBuffer_2_value;
    end
    if (sel) begin
      lineBuffer_4_grad_dir <= lineBuffer_3_grad_dir;
    end
    if (sel) begin
      lineBuffer_4_value <= lineBuffer_3_value;
    end
    if (sel) begin
      lineBuffer_5_grad_dir <= lineBuffer_4_grad_dir;
    end
    if (sel) begin
      lineBuffer_5_value <= lineBuffer_4_value;
    end
    if (sel) begin
      lineBuffer_6_grad_dir <= lineBuffer_5_grad_dir;
    end
    if (sel) begin
      lineBuffer_6_value <= lineBuffer_5_value;
    end
    if (sel) begin
      lineBuffer_7_grad_dir <= lineBuffer_6_grad_dir;
    end
    if (sel) begin
      lineBuffer_7_value <= lineBuffer_6_value;
    end
    if (sel) begin
      lineBuffer_8_grad_dir <= lineBuffer_7_grad_dir;
    end
    if (sel) begin
      lineBuffer_8_value <= lineBuffer_7_value;
    end
    if (sel) begin
      lineBuffer_9_grad_dir <= lineBuffer_8_grad_dir;
    end
    if (sel) begin
      lineBuffer_9_value <= lineBuffer_8_value;
    end
    if (sel) begin
      lineBuffer_10_grad_dir <= lineBuffer_9_grad_dir;
    end
    if (sel) begin
      lineBuffer_10_value <= lineBuffer_9_value;
    end
    if (sel) begin
      lineBuffer_11_grad_dir <= lineBuffer_10_grad_dir;
    end
    if (sel) begin
      lineBuffer_11_value <= lineBuffer_10_value;
    end
    if (sel) begin
      lineBuffer_12_grad_dir <= lineBuffer_11_grad_dir;
    end
    if (sel) begin
      lineBuffer_12_value <= lineBuffer_11_value;
    end
    if (sel) begin
      lineBuffer_13_grad_dir <= lineBuffer_12_grad_dir;
    end
    if (sel) begin
      lineBuffer_13_value <= lineBuffer_12_value;
    end
    if (sel) begin
      lineBuffer_14_grad_dir <= lineBuffer_13_grad_dir;
    end
    if (sel) begin
      lineBuffer_14_value <= lineBuffer_13_value;
    end
    if (sel) begin
      lineBuffer_15_grad_dir <= lineBuffer_14_grad_dir;
    end
    if (sel) begin
      lineBuffer_15_value <= lineBuffer_14_value;
    end
    if (sel) begin
      lineBuffer_16_grad_dir <= lineBuffer_15_grad_dir;
    end
    if (sel) begin
      lineBuffer_16_value <= lineBuffer_15_value;
    end
    if (sel) begin
      lineBuffer_17_grad_dir <= lineBuffer_16_grad_dir;
    end
    if (sel) begin
      lineBuffer_17_value <= lineBuffer_16_value;
    end
    if (sel) begin
      lineBuffer_18_grad_dir <= lineBuffer_17_grad_dir;
    end
    if (sel) begin
      lineBuffer_18_value <= lineBuffer_17_value;
    end
    if (sel) begin
      lineBuffer_19_grad_dir <= lineBuffer_18_grad_dir;
    end
    if (sel) begin
      lineBuffer_19_value <= lineBuffer_18_value;
    end
    if (sel) begin
      lineBuffer_20_grad_dir <= lineBuffer_19_grad_dir;
    end
    if (sel) begin
      lineBuffer_20_value <= lineBuffer_19_value;
    end
    if (sel) begin
      lineBuffer_21_grad_dir <= lineBuffer_20_grad_dir;
    end
    if (sel) begin
      lineBuffer_21_value <= lineBuffer_20_value;
    end
    if (sel) begin
      lineBuffer_22_grad_dir <= lineBuffer_21_grad_dir;
    end
    if (sel) begin
      lineBuffer_22_value <= lineBuffer_21_value;
    end
    if (sel) begin
      lineBuffer_23_grad_dir <= lineBuffer_22_grad_dir;
    end
    if (sel) begin
      lineBuffer_23_value <= lineBuffer_22_value;
    end
    if (sel) begin
      lineBuffer_24_grad_dir <= lineBuffer_23_grad_dir;
    end
    if (sel) begin
      lineBuffer_24_value <= lineBuffer_23_value;
    end
    if (sel) begin
      lineBuffer_25_grad_dir <= lineBuffer_24_grad_dir;
    end
    if (sel) begin
      lineBuffer_25_value <= lineBuffer_24_value;
    end
    if (sel) begin
      lineBuffer_26_grad_dir <= lineBuffer_25_grad_dir;
    end
    if (sel) begin
      lineBuffer_26_value <= lineBuffer_25_value;
    end
    if (sel) begin
      lineBuffer_27_grad_dir <= lineBuffer_26_grad_dir;
    end
    if (sel) begin
      lineBuffer_27_value <= lineBuffer_26_value;
    end
    if (sel) begin
      lineBuffer_28_grad_dir <= lineBuffer_27_grad_dir;
    end
    if (sel) begin
      lineBuffer_28_value <= lineBuffer_27_value;
    end
    if (sel) begin
      lineBuffer_29_grad_dir <= lineBuffer_28_grad_dir;
    end
    if (sel) begin
      lineBuffer_29_value <= lineBuffer_28_value;
    end
    if (sel) begin
      lineBuffer_30_grad_dir <= lineBuffer_29_grad_dir;
    end
    if (sel) begin
      lineBuffer_30_value <= lineBuffer_29_value;
    end
    if (sel) begin
      lineBuffer_31_grad_dir <= lineBuffer_30_grad_dir;
    end
    if (sel) begin
      lineBuffer_31_value <= lineBuffer_30_value;
    end
    if (sel) begin
      lineBuffer_32_grad_dir <= lineBuffer_31_grad_dir;
    end
    if (sel) begin
      lineBuffer_32_value <= lineBuffer_31_value;
    end
    if (sel) begin
      lineBuffer_33_grad_dir <= lineBuffer_32_grad_dir;
    end
    if (sel) begin
      lineBuffer_33_value <= lineBuffer_32_value;
    end
    if (sel) begin
      lineBuffer_34_grad_dir <= lineBuffer_33_grad_dir;
    end
    if (sel) begin
      lineBuffer_34_value <= lineBuffer_33_value;
    end
    if (sel) begin
      lineBuffer_35_grad_dir <= lineBuffer_34_grad_dir;
    end
    if (sel) begin
      lineBuffer_35_value <= lineBuffer_34_value;
    end
    if (sel) begin
      lineBuffer_36_grad_dir <= lineBuffer_35_grad_dir;
    end
    if (sel) begin
      lineBuffer_36_value <= lineBuffer_35_value;
    end
    if (sel) begin
      lineBuffer_37_grad_dir <= lineBuffer_36_grad_dir;
    end
    if (sel) begin
      lineBuffer_37_value <= lineBuffer_36_value;
    end
    if (sel) begin
      lineBuffer_38_grad_dir <= lineBuffer_37_grad_dir;
    end
    if (sel) begin
      lineBuffer_38_value <= lineBuffer_37_value;
    end
    if (sel) begin
      lineBuffer_39_grad_dir <= lineBuffer_38_grad_dir;
    end
    if (sel) begin
      lineBuffer_39_value <= lineBuffer_38_value;
    end
    if (sel) begin
      lineBuffer_40_grad_dir <= lineBuffer_39_grad_dir;
    end
    if (sel) begin
      lineBuffer_40_value <= lineBuffer_39_value;
    end
    if (sel) begin
      lineBuffer_41_grad_dir <= lineBuffer_40_grad_dir;
    end
    if (sel) begin
      lineBuffer_41_value <= lineBuffer_40_value;
    end
    if (sel) begin
      lineBuffer_42_grad_dir <= lineBuffer_41_grad_dir;
    end
    if (sel) begin
      lineBuffer_42_value <= lineBuffer_41_value;
    end
    if (sel) begin
      lineBuffer_43_grad_dir <= lineBuffer_42_grad_dir;
    end
    if (sel) begin
      lineBuffer_43_value <= lineBuffer_42_value;
    end
    if (sel) begin
      lineBuffer_44_grad_dir <= lineBuffer_43_grad_dir;
    end
    if (sel) begin
      lineBuffer_44_value <= lineBuffer_43_value;
    end
    if (sel) begin
      lineBuffer_45_grad_dir <= lineBuffer_44_grad_dir;
    end
    if (sel) begin
      lineBuffer_45_value <= lineBuffer_44_value;
    end
    if (sel) begin
      lineBuffer_46_grad_dir <= lineBuffer_45_grad_dir;
    end
    if (sel) begin
      lineBuffer_46_value <= lineBuffer_45_value;
    end
    if (sel) begin
      lineBuffer_47_grad_dir <= lineBuffer_46_grad_dir;
    end
    if (sel) begin
      lineBuffer_47_value <= lineBuffer_46_value;
    end
    if (sel) begin
      lineBuffer_48_grad_dir <= lineBuffer_47_grad_dir;
    end
    if (sel) begin
      lineBuffer_48_value <= lineBuffer_47_value;
    end
    if (sel) begin
      lineBuffer_49_grad_dir <= lineBuffer_48_grad_dir;
    end
    if (sel) begin
      lineBuffer_49_value <= lineBuffer_48_value;
    end
    if (sel) begin
      lineBuffer_50_grad_dir <= lineBuffer_49_grad_dir;
    end
    if (sel) begin
      lineBuffer_50_value <= lineBuffer_49_value;
    end
    if (sel) begin
      lineBuffer_51_grad_dir <= lineBuffer_50_grad_dir;
    end
    if (sel) begin
      lineBuffer_51_value <= lineBuffer_50_value;
    end
    if (sel) begin
      lineBuffer_52_grad_dir <= lineBuffer_51_grad_dir;
    end
    if (sel) begin
      lineBuffer_52_value <= lineBuffer_51_value;
    end
    if (sel) begin
      lineBuffer_53_grad_dir <= lineBuffer_52_grad_dir;
    end
    if (sel) begin
      lineBuffer_53_value <= lineBuffer_52_value;
    end
    if (sel) begin
      lineBuffer_54_grad_dir <= lineBuffer_53_grad_dir;
    end
    if (sel) begin
      lineBuffer_54_value <= lineBuffer_53_value;
    end
    if (sel) begin
      lineBuffer_55_grad_dir <= lineBuffer_54_grad_dir;
    end
    if (sel) begin
      lineBuffer_55_value <= lineBuffer_54_value;
    end
    if (sel) begin
      lineBuffer_56_grad_dir <= lineBuffer_55_grad_dir;
    end
    if (sel) begin
      lineBuffer_56_value <= lineBuffer_55_value;
    end
    if (sel) begin
      lineBuffer_57_grad_dir <= lineBuffer_56_grad_dir;
    end
    if (sel) begin
      lineBuffer_57_value <= lineBuffer_56_value;
    end
    if (sel) begin
      lineBuffer_58_grad_dir <= lineBuffer_57_grad_dir;
    end
    if (sel) begin
      lineBuffer_58_value <= lineBuffer_57_value;
    end
    if (sel) begin
      lineBuffer_59_grad_dir <= lineBuffer_58_grad_dir;
    end
    if (sel) begin
      lineBuffer_59_value <= lineBuffer_58_value;
    end
    if (sel) begin
      lineBuffer_60_grad_dir <= lineBuffer_59_grad_dir;
    end
    if (sel) begin
      lineBuffer_60_value <= lineBuffer_59_value;
    end
    if (sel) begin
      lineBuffer_61_grad_dir <= lineBuffer_60_grad_dir;
    end
    if (sel) begin
      lineBuffer_61_value <= lineBuffer_60_value;
    end
    if (sel) begin
      lineBuffer_62_grad_dir <= lineBuffer_61_grad_dir;
    end
    if (sel) begin
      lineBuffer_62_value <= lineBuffer_61_value;
    end
    if (sel) begin
      lineBuffer_63_grad_dir <= lineBuffer_62_grad_dir;
    end
    if (sel) begin
      lineBuffer_63_value <= lineBuffer_62_value;
    end
    if (sel) begin
      lineBuffer_64_grad_dir <= lineBuffer_63_grad_dir;
    end
    if (sel) begin
      lineBuffer_64_value <= lineBuffer_63_value;
    end
    if (sel) begin
      lineBuffer_65_grad_dir <= lineBuffer_64_grad_dir;
    end
    if (sel) begin
      lineBuffer_65_value <= lineBuffer_64_value;
    end
    if (sel) begin
      lineBuffer_66_grad_dir <= lineBuffer_65_grad_dir;
    end
    if (sel) begin
      lineBuffer_66_value <= lineBuffer_65_value;
    end
    if (sel) begin
      lineBuffer_67_grad_dir <= lineBuffer_66_grad_dir;
    end
    if (sel) begin
      lineBuffer_67_value <= lineBuffer_66_value;
    end
    if (sel) begin
      lineBuffer_68_grad_dir <= lineBuffer_67_grad_dir;
    end
    if (sel) begin
      lineBuffer_68_value <= lineBuffer_67_value;
    end
    if (sel) begin
      lineBuffer_69_grad_dir <= lineBuffer_68_grad_dir;
    end
    if (sel) begin
      lineBuffer_69_value <= lineBuffer_68_value;
    end
    if (sel) begin
      lineBuffer_70_grad_dir <= lineBuffer_69_grad_dir;
    end
    if (sel) begin
      lineBuffer_70_value <= lineBuffer_69_value;
    end
    if (sel) begin
      lineBuffer_71_grad_dir <= lineBuffer_70_grad_dir;
    end
    if (sel) begin
      lineBuffer_71_value <= lineBuffer_70_value;
    end
    if (sel) begin
      lineBuffer_72_grad_dir <= lineBuffer_71_grad_dir;
    end
    if (sel) begin
      lineBuffer_72_value <= lineBuffer_71_value;
    end
    if (sel) begin
      lineBuffer_73_grad_dir <= lineBuffer_72_grad_dir;
    end
    if (sel) begin
      lineBuffer_73_value <= lineBuffer_72_value;
    end
    if (sel) begin
      lineBuffer_74_grad_dir <= lineBuffer_73_grad_dir;
    end
    if (sel) begin
      lineBuffer_74_value <= lineBuffer_73_value;
    end
    if (sel) begin
      lineBuffer_75_grad_dir <= lineBuffer_74_grad_dir;
    end
    if (sel) begin
      lineBuffer_75_value <= lineBuffer_74_value;
    end
    if (sel) begin
      lineBuffer_76_grad_dir <= lineBuffer_75_grad_dir;
    end
    if (sel) begin
      lineBuffer_76_value <= lineBuffer_75_value;
    end
    if (sel) begin
      lineBuffer_77_grad_dir <= lineBuffer_76_grad_dir;
    end
    if (sel) begin
      lineBuffer_77_value <= lineBuffer_76_value;
    end
    if (sel) begin
      lineBuffer_78_grad_dir <= lineBuffer_77_grad_dir;
    end
    if (sel) begin
      lineBuffer_78_value <= lineBuffer_77_value;
    end
    if (sel) begin
      lineBuffer_79_grad_dir <= lineBuffer_78_grad_dir;
    end
    if (sel) begin
      lineBuffer_79_value <= lineBuffer_78_value;
    end
    if (sel) begin
      lineBuffer_80_grad_dir <= lineBuffer_79_grad_dir;
    end
    if (sel) begin
      lineBuffer_80_value <= lineBuffer_79_value;
    end
    if (sel) begin
      lineBuffer_81_grad_dir <= lineBuffer_80_grad_dir;
    end
    if (sel) begin
      lineBuffer_81_value <= lineBuffer_80_value;
    end
    if (sel) begin
      lineBuffer_82_grad_dir <= lineBuffer_81_grad_dir;
    end
    if (sel) begin
      lineBuffer_82_value <= lineBuffer_81_value;
    end
    if (sel) begin
      lineBuffer_83_grad_dir <= lineBuffer_82_grad_dir;
    end
    if (sel) begin
      lineBuffer_83_value <= lineBuffer_82_value;
    end
    if (sel) begin
      lineBuffer_84_grad_dir <= lineBuffer_83_grad_dir;
    end
    if (sel) begin
      lineBuffer_84_value <= lineBuffer_83_value;
    end
    if (sel) begin
      lineBuffer_85_grad_dir <= lineBuffer_84_grad_dir;
    end
    if (sel) begin
      lineBuffer_85_value <= lineBuffer_84_value;
    end
    if (sel) begin
      lineBuffer_86_grad_dir <= lineBuffer_85_grad_dir;
    end
    if (sel) begin
      lineBuffer_86_value <= lineBuffer_85_value;
    end
    if (sel) begin
      lineBuffer_87_grad_dir <= lineBuffer_86_grad_dir;
    end
    if (sel) begin
      lineBuffer_87_value <= lineBuffer_86_value;
    end
    if (sel) begin
      lineBuffer_88_grad_dir <= lineBuffer_87_grad_dir;
    end
    if (sel) begin
      lineBuffer_88_value <= lineBuffer_87_value;
    end
    if (sel) begin
      lineBuffer_89_grad_dir <= lineBuffer_88_grad_dir;
    end
    if (sel) begin
      lineBuffer_89_value <= lineBuffer_88_value;
    end
    if (sel) begin
      lineBuffer_90_grad_dir <= lineBuffer_89_grad_dir;
    end
    if (sel) begin
      lineBuffer_90_value <= lineBuffer_89_value;
    end
    if (sel) begin
      lineBuffer_91_grad_dir <= lineBuffer_90_grad_dir;
    end
    if (sel) begin
      lineBuffer_91_value <= lineBuffer_90_value;
    end
    if (sel) begin
      lineBuffer_92_grad_dir <= lineBuffer_91_grad_dir;
    end
    if (sel) begin
      lineBuffer_92_value <= lineBuffer_91_value;
    end
    if (sel) begin
      lineBuffer_93_grad_dir <= lineBuffer_92_grad_dir;
    end
    if (sel) begin
      lineBuffer_93_value <= lineBuffer_92_value;
    end
    if (sel) begin
      lineBuffer_94_grad_dir <= lineBuffer_93_grad_dir;
    end
    if (sel) begin
      lineBuffer_94_value <= lineBuffer_93_value;
    end
    if (sel) begin
      lineBuffer_95_grad_dir <= lineBuffer_94_grad_dir;
    end
    if (sel) begin
      lineBuffer_95_value <= lineBuffer_94_value;
    end
    if (sel) begin
      lineBuffer_96_grad_dir <= lineBuffer_95_grad_dir;
    end
    if (sel) begin
      lineBuffer_96_value <= lineBuffer_95_value;
    end
    if (sel) begin
      lineBuffer_97_grad_dir <= lineBuffer_96_grad_dir;
    end
    if (sel) begin
      lineBuffer_97_value <= lineBuffer_96_value;
    end
    if (sel) begin
      lineBuffer_98_grad_dir <= lineBuffer_97_grad_dir;
    end
    if (sel) begin
      lineBuffer_98_value <= lineBuffer_97_value;
    end
    if (sel) begin
      lineBuffer_99_grad_dir <= lineBuffer_98_grad_dir;
    end
    if (sel) begin
      lineBuffer_99_value <= lineBuffer_98_value;
    end
    if (sel) begin
      lineBuffer_100_grad_dir <= lineBuffer_99_grad_dir;
    end
    if (sel) begin
      lineBuffer_100_value <= lineBuffer_99_value;
    end
    if (sel) begin
      lineBuffer_101_grad_dir <= lineBuffer_100_grad_dir;
    end
    if (sel) begin
      lineBuffer_101_value <= lineBuffer_100_value;
    end
    if (sel) begin
      lineBuffer_102_grad_dir <= lineBuffer_101_grad_dir;
    end
    if (sel) begin
      lineBuffer_102_value <= lineBuffer_101_value;
    end
    if (sel) begin
      lineBuffer_103_grad_dir <= lineBuffer_102_grad_dir;
    end
    if (sel) begin
      lineBuffer_103_value <= lineBuffer_102_value;
    end
    if (sel) begin
      lineBuffer_104_grad_dir <= lineBuffer_103_grad_dir;
    end
    if (sel) begin
      lineBuffer_104_value <= lineBuffer_103_value;
    end
    if (sel) begin
      lineBuffer_105_grad_dir <= lineBuffer_104_grad_dir;
    end
    if (sel) begin
      lineBuffer_105_value <= lineBuffer_104_value;
    end
    if (sel) begin
      lineBuffer_106_grad_dir <= lineBuffer_105_grad_dir;
    end
    if (sel) begin
      lineBuffer_106_value <= lineBuffer_105_value;
    end
    if (sel) begin
      lineBuffer_107_grad_dir <= lineBuffer_106_grad_dir;
    end
    if (sel) begin
      lineBuffer_107_value <= lineBuffer_106_value;
    end
    if (sel) begin
      lineBuffer_108_grad_dir <= lineBuffer_107_grad_dir;
    end
    if (sel) begin
      lineBuffer_108_value <= lineBuffer_107_value;
    end
    if (sel) begin
      lineBuffer_109_grad_dir <= lineBuffer_108_grad_dir;
    end
    if (sel) begin
      lineBuffer_109_value <= lineBuffer_108_value;
    end
    if (sel) begin
      lineBuffer_110_grad_dir <= lineBuffer_109_grad_dir;
    end
    if (sel) begin
      lineBuffer_110_value <= lineBuffer_109_value;
    end
    if (sel) begin
      lineBuffer_111_grad_dir <= lineBuffer_110_grad_dir;
    end
    if (sel) begin
      lineBuffer_111_value <= lineBuffer_110_value;
    end
    if (sel) begin
      lineBuffer_112_grad_dir <= lineBuffer_111_grad_dir;
    end
    if (sel) begin
      lineBuffer_112_value <= lineBuffer_111_value;
    end
    if (sel) begin
      lineBuffer_113_grad_dir <= lineBuffer_112_grad_dir;
    end
    if (sel) begin
      lineBuffer_113_value <= lineBuffer_112_value;
    end
    if (sel) begin
      lineBuffer_114_grad_dir <= lineBuffer_113_grad_dir;
    end
    if (sel) begin
      lineBuffer_114_value <= lineBuffer_113_value;
    end
    if (sel) begin
      lineBuffer_115_grad_dir <= lineBuffer_114_grad_dir;
    end
    if (sel) begin
      lineBuffer_115_value <= lineBuffer_114_value;
    end
    if (sel) begin
      lineBuffer_116_grad_dir <= lineBuffer_115_grad_dir;
    end
    if (sel) begin
      lineBuffer_116_value <= lineBuffer_115_value;
    end
    if (sel) begin
      lineBuffer_117_grad_dir <= lineBuffer_116_grad_dir;
    end
    if (sel) begin
      lineBuffer_117_value <= lineBuffer_116_value;
    end
    if (sel) begin
      lineBuffer_118_grad_dir <= lineBuffer_117_grad_dir;
    end
    if (sel) begin
      lineBuffer_118_value <= lineBuffer_117_value;
    end
    if (sel) begin
      lineBuffer_119_grad_dir <= lineBuffer_118_grad_dir;
    end
    if (sel) begin
      lineBuffer_119_value <= lineBuffer_118_value;
    end
    if (sel) begin
      lineBuffer_120_grad_dir <= lineBuffer_119_grad_dir;
    end
    if (sel) begin
      lineBuffer_120_value <= lineBuffer_119_value;
    end
    if (sel) begin
      lineBuffer_121_grad_dir <= lineBuffer_120_grad_dir;
    end
    if (sel) begin
      lineBuffer_121_value <= lineBuffer_120_value;
    end
    if (sel) begin
      lineBuffer_122_grad_dir <= lineBuffer_121_grad_dir;
    end
    if (sel) begin
      lineBuffer_122_value <= lineBuffer_121_value;
    end
    if (sel) begin
      lineBuffer_123_grad_dir <= lineBuffer_122_grad_dir;
    end
    if (sel) begin
      lineBuffer_123_value <= lineBuffer_122_value;
    end
    if (sel) begin
      lineBuffer_124_grad_dir <= lineBuffer_123_grad_dir;
    end
    if (sel) begin
      lineBuffer_124_value <= lineBuffer_123_value;
    end
    if (sel) begin
      lineBuffer_125_grad_dir <= lineBuffer_124_grad_dir;
    end
    if (sel) begin
      lineBuffer_125_value <= lineBuffer_124_value;
    end
    if (sel) begin
      lineBuffer_126_grad_dir <= lineBuffer_125_grad_dir;
    end
    if (sel) begin
      lineBuffer_126_value <= lineBuffer_125_value;
    end
    if (sel) begin
      lineBuffer_127_grad_dir <= lineBuffer_126_grad_dir;
    end
    if (sel) begin
      lineBuffer_127_value <= lineBuffer_126_value;
    end
    if (sel) begin
      lineBuffer_128_grad_dir <= lineBuffer_127_grad_dir;
    end
    if (sel) begin
      lineBuffer_128_value <= lineBuffer_127_value;
    end
    if (sel) begin
      lineBuffer_129_grad_dir <= lineBuffer_128_grad_dir;
    end
    if (sel) begin
      lineBuffer_129_value <= lineBuffer_128_value;
    end
    if (sel) begin
      lineBuffer_130_grad_dir <= lineBuffer_129_grad_dir;
    end
    if (sel) begin
      lineBuffer_130_value <= lineBuffer_129_value;
    end
    if (sel) begin
      lineBuffer_131_grad_dir <= lineBuffer_130_grad_dir;
    end
    if (sel) begin
      lineBuffer_131_value <= lineBuffer_130_value;
    end
    if (sel) begin
      lineBuffer_132_grad_dir <= lineBuffer_131_grad_dir;
    end
    if (sel) begin
      lineBuffer_132_value <= lineBuffer_131_value;
    end
    if (sel) begin
      lineBuffer_133_grad_dir <= lineBuffer_132_grad_dir;
    end
    if (sel) begin
      lineBuffer_133_value <= lineBuffer_132_value;
    end
    if (sel) begin
      lineBuffer_134_grad_dir <= lineBuffer_133_grad_dir;
    end
    if (sel) begin
      lineBuffer_134_value <= lineBuffer_133_value;
    end
    if (sel) begin
      lineBuffer_135_grad_dir <= lineBuffer_134_grad_dir;
    end
    if (sel) begin
      lineBuffer_135_value <= lineBuffer_134_value;
    end
    if (sel) begin
      lineBuffer_136_grad_dir <= lineBuffer_135_grad_dir;
    end
    if (sel) begin
      lineBuffer_136_value <= lineBuffer_135_value;
    end
    if (sel) begin
      lineBuffer_137_grad_dir <= lineBuffer_136_grad_dir;
    end
    if (sel) begin
      lineBuffer_137_value <= lineBuffer_136_value;
    end
    if (sel) begin
      lineBuffer_138_grad_dir <= lineBuffer_137_grad_dir;
    end
    if (sel) begin
      lineBuffer_138_value <= lineBuffer_137_value;
    end
    if (sel) begin
      lineBuffer_139_grad_dir <= lineBuffer_138_grad_dir;
    end
    if (sel) begin
      lineBuffer_139_value <= lineBuffer_138_value;
    end
    if (sel) begin
      lineBuffer_140_grad_dir <= lineBuffer_139_grad_dir;
    end
    if (sel) begin
      lineBuffer_140_value <= lineBuffer_139_value;
    end
    if (sel) begin
      lineBuffer_141_grad_dir <= lineBuffer_140_grad_dir;
    end
    if (sel) begin
      lineBuffer_141_value <= lineBuffer_140_value;
    end
    if (sel) begin
      lineBuffer_142_grad_dir <= lineBuffer_141_grad_dir;
    end
    if (sel) begin
      lineBuffer_142_value <= lineBuffer_141_value;
    end
    if (sel) begin
      lineBuffer_143_grad_dir <= lineBuffer_142_grad_dir;
    end
    if (sel) begin
      lineBuffer_143_value <= lineBuffer_142_value;
    end
    if (sel) begin
      lineBuffer_144_grad_dir <= lineBuffer_143_grad_dir;
    end
    if (sel) begin
      lineBuffer_144_value <= lineBuffer_143_value;
    end
    if (sel) begin
      lineBuffer_145_grad_dir <= lineBuffer_144_grad_dir;
    end
    if (sel) begin
      lineBuffer_145_value <= lineBuffer_144_value;
    end
    if (sel) begin
      lineBuffer_146_grad_dir <= lineBuffer_145_grad_dir;
    end
    if (sel) begin
      lineBuffer_146_value <= lineBuffer_145_value;
    end
    if (sel) begin
      lineBuffer_147_grad_dir <= lineBuffer_146_grad_dir;
    end
    if (sel) begin
      lineBuffer_147_value <= lineBuffer_146_value;
    end
    if (sel) begin
      lineBuffer_148_grad_dir <= lineBuffer_147_grad_dir;
    end
    if (sel) begin
      lineBuffer_148_value <= lineBuffer_147_value;
    end
    if (sel) begin
      lineBuffer_149_grad_dir <= lineBuffer_148_grad_dir;
    end
    if (sel) begin
      lineBuffer_149_value <= lineBuffer_148_value;
    end
    if (sel) begin
      lineBuffer_150_grad_dir <= lineBuffer_149_grad_dir;
    end
    if (sel) begin
      lineBuffer_150_value <= lineBuffer_149_value;
    end
    if (sel) begin
      lineBuffer_151_grad_dir <= lineBuffer_150_grad_dir;
    end
    if (sel) begin
      lineBuffer_151_value <= lineBuffer_150_value;
    end
    if (sel) begin
      lineBuffer_152_grad_dir <= lineBuffer_151_grad_dir;
    end
    if (sel) begin
      lineBuffer_152_value <= lineBuffer_151_value;
    end
    if (sel) begin
      lineBuffer_153_grad_dir <= lineBuffer_152_grad_dir;
    end
    if (sel) begin
      lineBuffer_153_value <= lineBuffer_152_value;
    end
    if (sel) begin
      lineBuffer_154_grad_dir <= lineBuffer_153_grad_dir;
    end
    if (sel) begin
      lineBuffer_154_value <= lineBuffer_153_value;
    end
    if (sel) begin
      lineBuffer_155_grad_dir <= lineBuffer_154_grad_dir;
    end
    if (sel) begin
      lineBuffer_155_value <= lineBuffer_154_value;
    end
    if (sel) begin
      lineBuffer_156_grad_dir <= lineBuffer_155_grad_dir;
    end
    if (sel) begin
      lineBuffer_156_value <= lineBuffer_155_value;
    end
    if (sel) begin
      lineBuffer_157_grad_dir <= lineBuffer_156_grad_dir;
    end
    if (sel) begin
      lineBuffer_157_value <= lineBuffer_156_value;
    end
    if (sel) begin
      lineBuffer_158_grad_dir <= lineBuffer_157_grad_dir;
    end
    if (sel) begin
      lineBuffer_158_value <= lineBuffer_157_value;
    end
    if (sel) begin
      lineBuffer_159_grad_dir <= lineBuffer_158_grad_dir;
    end
    if (sel) begin
      lineBuffer_159_value <= lineBuffer_158_value;
    end
    if (sel) begin
      lineBuffer_160_grad_dir <= lineBuffer_159_grad_dir;
    end
    if (sel) begin
      lineBuffer_160_value <= lineBuffer_159_value;
    end
    if (sel) begin
      lineBuffer_161_grad_dir <= lineBuffer_160_grad_dir;
    end
    if (sel) begin
      lineBuffer_161_value <= lineBuffer_160_value;
    end
    if (sel) begin
      lineBuffer_162_grad_dir <= lineBuffer_161_grad_dir;
    end
    if (sel) begin
      lineBuffer_162_value <= lineBuffer_161_value;
    end
    if (sel) begin
      lineBuffer_163_grad_dir <= lineBuffer_162_grad_dir;
    end
    if (sel) begin
      lineBuffer_163_value <= lineBuffer_162_value;
    end
    if (sel) begin
      lineBuffer_164_grad_dir <= lineBuffer_163_grad_dir;
    end
    if (sel) begin
      lineBuffer_164_value <= lineBuffer_163_value;
    end
    if (sel) begin
      lineBuffer_165_grad_dir <= lineBuffer_164_grad_dir;
    end
    if (sel) begin
      lineBuffer_165_value <= lineBuffer_164_value;
    end
    if (sel) begin
      lineBuffer_166_grad_dir <= lineBuffer_165_grad_dir;
    end
    if (sel) begin
      lineBuffer_166_value <= lineBuffer_165_value;
    end
    if (sel) begin
      lineBuffer_167_grad_dir <= lineBuffer_166_grad_dir;
    end
    if (sel) begin
      lineBuffer_167_value <= lineBuffer_166_value;
    end
    if (sel) begin
      lineBuffer_168_grad_dir <= lineBuffer_167_grad_dir;
    end
    if (sel) begin
      lineBuffer_168_value <= lineBuffer_167_value;
    end
    if (sel) begin
      lineBuffer_169_grad_dir <= lineBuffer_168_grad_dir;
    end
    if (sel) begin
      lineBuffer_169_value <= lineBuffer_168_value;
    end
    if (sel) begin
      lineBuffer_170_grad_dir <= lineBuffer_169_grad_dir;
    end
    if (sel) begin
      lineBuffer_170_value <= lineBuffer_169_value;
    end
    if (sel) begin
      lineBuffer_171_grad_dir <= lineBuffer_170_grad_dir;
    end
    if (sel) begin
      lineBuffer_171_value <= lineBuffer_170_value;
    end
    if (sel) begin
      lineBuffer_172_grad_dir <= lineBuffer_171_grad_dir;
    end
    if (sel) begin
      lineBuffer_172_value <= lineBuffer_171_value;
    end
    if (sel) begin
      lineBuffer_173_grad_dir <= lineBuffer_172_grad_dir;
    end
    if (sel) begin
      lineBuffer_173_value <= lineBuffer_172_value;
    end
    if (sel) begin
      lineBuffer_174_grad_dir <= lineBuffer_173_grad_dir;
    end
    if (sel) begin
      lineBuffer_174_value <= lineBuffer_173_value;
    end
    if (sel) begin
      lineBuffer_175_grad_dir <= lineBuffer_174_grad_dir;
    end
    if (sel) begin
      lineBuffer_175_value <= lineBuffer_174_value;
    end
    if (sel) begin
      lineBuffer_176_grad_dir <= lineBuffer_175_grad_dir;
    end
    if (sel) begin
      lineBuffer_176_value <= lineBuffer_175_value;
    end
    if (sel) begin
      lineBuffer_177_grad_dir <= lineBuffer_176_grad_dir;
    end
    if (sel) begin
      lineBuffer_177_value <= lineBuffer_176_value;
    end
    if (sel) begin
      lineBuffer_178_grad_dir <= lineBuffer_177_grad_dir;
    end
    if (sel) begin
      lineBuffer_178_value <= lineBuffer_177_value;
    end
    if (sel) begin
      lineBuffer_179_grad_dir <= lineBuffer_178_grad_dir;
    end
    if (sel) begin
      lineBuffer_179_value <= lineBuffer_178_value;
    end
    if (sel) begin
      lineBuffer_180_grad_dir <= lineBuffer_179_grad_dir;
    end
    if (sel) begin
      lineBuffer_180_value <= lineBuffer_179_value;
    end
    if (sel) begin
      lineBuffer_181_grad_dir <= lineBuffer_180_grad_dir;
    end
    if (sel) begin
      lineBuffer_181_value <= lineBuffer_180_value;
    end
    if (sel) begin
      lineBuffer_182_grad_dir <= lineBuffer_181_grad_dir;
    end
    if (sel) begin
      lineBuffer_182_value <= lineBuffer_181_value;
    end
    if (sel) begin
      lineBuffer_183_grad_dir <= lineBuffer_182_grad_dir;
    end
    if (sel) begin
      lineBuffer_183_value <= lineBuffer_182_value;
    end
    if (sel) begin
      lineBuffer_184_grad_dir <= lineBuffer_183_grad_dir;
    end
    if (sel) begin
      lineBuffer_184_value <= lineBuffer_183_value;
    end
    if (sel) begin
      lineBuffer_185_grad_dir <= lineBuffer_184_grad_dir;
    end
    if (sel) begin
      lineBuffer_185_value <= lineBuffer_184_value;
    end
    if (sel) begin
      lineBuffer_186_grad_dir <= lineBuffer_185_grad_dir;
    end
    if (sel) begin
      lineBuffer_186_value <= lineBuffer_185_value;
    end
    if (sel) begin
      lineBuffer_187_grad_dir <= lineBuffer_186_grad_dir;
    end
    if (sel) begin
      lineBuffer_187_value <= lineBuffer_186_value;
    end
    if (sel) begin
      lineBuffer_188_grad_dir <= lineBuffer_187_grad_dir;
    end
    if (sel) begin
      lineBuffer_188_value <= lineBuffer_187_value;
    end
    if (sel) begin
      lineBuffer_189_grad_dir <= lineBuffer_188_grad_dir;
    end
    if (sel) begin
      lineBuffer_189_value <= lineBuffer_188_value;
    end
    if (sel) begin
      lineBuffer_190_grad_dir <= lineBuffer_189_grad_dir;
    end
    if (sel) begin
      lineBuffer_190_value <= lineBuffer_189_value;
    end
    if (sel) begin
      lineBuffer_191_grad_dir <= lineBuffer_190_grad_dir;
    end
    if (sel) begin
      lineBuffer_191_value <= lineBuffer_190_value;
    end
    if (sel) begin
      lineBuffer_192_grad_dir <= lineBuffer_191_grad_dir;
    end
    if (sel) begin
      lineBuffer_192_value <= lineBuffer_191_value;
    end
    if (sel) begin
      lineBuffer_193_grad_dir <= lineBuffer_192_grad_dir;
    end
    if (sel) begin
      lineBuffer_193_value <= lineBuffer_192_value;
    end
    if (sel) begin
      lineBuffer_194_grad_dir <= lineBuffer_193_grad_dir;
    end
    if (sel) begin
      lineBuffer_194_value <= lineBuffer_193_value;
    end
    if (sel) begin
      lineBuffer_195_grad_dir <= lineBuffer_194_grad_dir;
    end
    if (sel) begin
      lineBuffer_195_value <= lineBuffer_194_value;
    end
    if (sel) begin
      lineBuffer_196_grad_dir <= lineBuffer_195_grad_dir;
    end
    if (sel) begin
      lineBuffer_196_value <= lineBuffer_195_value;
    end
    if (sel) begin
      lineBuffer_197_grad_dir <= lineBuffer_196_grad_dir;
    end
    if (sel) begin
      lineBuffer_197_value <= lineBuffer_196_value;
    end
    if (sel) begin
      lineBuffer_198_grad_dir <= lineBuffer_197_grad_dir;
    end
    if (sel) begin
      lineBuffer_198_value <= lineBuffer_197_value;
    end
    if (sel) begin
      lineBuffer_199_grad_dir <= lineBuffer_198_grad_dir;
    end
    if (sel) begin
      lineBuffer_199_value <= lineBuffer_198_value;
    end
    if (sel) begin
      lineBuffer_200_grad_dir <= lineBuffer_199_grad_dir;
    end
    if (sel) begin
      lineBuffer_200_value <= lineBuffer_199_value;
    end
    if (sel) begin
      lineBuffer_201_grad_dir <= lineBuffer_200_grad_dir;
    end
    if (sel) begin
      lineBuffer_201_value <= lineBuffer_200_value;
    end
    if (sel) begin
      lineBuffer_202_grad_dir <= lineBuffer_201_grad_dir;
    end
    if (sel) begin
      lineBuffer_202_value <= lineBuffer_201_value;
    end
    if (sel) begin
      lineBuffer_203_grad_dir <= lineBuffer_202_grad_dir;
    end
    if (sel) begin
      lineBuffer_203_value <= lineBuffer_202_value;
    end
    if (sel) begin
      lineBuffer_204_grad_dir <= lineBuffer_203_grad_dir;
    end
    if (sel) begin
      lineBuffer_204_value <= lineBuffer_203_value;
    end
    if (sel) begin
      lineBuffer_205_grad_dir <= lineBuffer_204_grad_dir;
    end
    if (sel) begin
      lineBuffer_205_value <= lineBuffer_204_value;
    end
    if (sel) begin
      lineBuffer_206_grad_dir <= lineBuffer_205_grad_dir;
    end
    if (sel) begin
      lineBuffer_206_value <= lineBuffer_205_value;
    end
    if (sel) begin
      lineBuffer_207_grad_dir <= lineBuffer_206_grad_dir;
    end
    if (sel) begin
      lineBuffer_207_value <= lineBuffer_206_value;
    end
    if (sel) begin
      lineBuffer_208_grad_dir <= lineBuffer_207_grad_dir;
    end
    if (sel) begin
      lineBuffer_208_value <= lineBuffer_207_value;
    end
    if (sel) begin
      lineBuffer_209_grad_dir <= lineBuffer_208_grad_dir;
    end
    if (sel) begin
      lineBuffer_209_value <= lineBuffer_208_value;
    end
    if (sel) begin
      lineBuffer_210_grad_dir <= lineBuffer_209_grad_dir;
    end
    if (sel) begin
      lineBuffer_210_value <= lineBuffer_209_value;
    end
    if (sel) begin
      lineBuffer_211_grad_dir <= lineBuffer_210_grad_dir;
    end
    if (sel) begin
      lineBuffer_211_value <= lineBuffer_210_value;
    end
    if (sel) begin
      lineBuffer_212_grad_dir <= lineBuffer_211_grad_dir;
    end
    if (sel) begin
      lineBuffer_212_value <= lineBuffer_211_value;
    end
    if (sel) begin
      lineBuffer_213_grad_dir <= lineBuffer_212_grad_dir;
    end
    if (sel) begin
      lineBuffer_213_value <= lineBuffer_212_value;
    end
    if (sel) begin
      lineBuffer_214_grad_dir <= lineBuffer_213_grad_dir;
    end
    if (sel) begin
      lineBuffer_214_value <= lineBuffer_213_value;
    end
    if (sel) begin
      lineBuffer_215_grad_dir <= lineBuffer_214_grad_dir;
    end
    if (sel) begin
      lineBuffer_215_value <= lineBuffer_214_value;
    end
    if (sel) begin
      lineBuffer_216_grad_dir <= lineBuffer_215_grad_dir;
    end
    if (sel) begin
      lineBuffer_216_value <= lineBuffer_215_value;
    end
    if (sel) begin
      lineBuffer_217_grad_dir <= lineBuffer_216_grad_dir;
    end
    if (sel) begin
      lineBuffer_217_value <= lineBuffer_216_value;
    end
    if (sel) begin
      lineBuffer_218_grad_dir <= lineBuffer_217_grad_dir;
    end
    if (sel) begin
      lineBuffer_218_value <= lineBuffer_217_value;
    end
    if (sel) begin
      lineBuffer_219_grad_dir <= lineBuffer_218_grad_dir;
    end
    if (sel) begin
      lineBuffer_219_value <= lineBuffer_218_value;
    end
    if (sel) begin
      lineBuffer_220_grad_dir <= lineBuffer_219_grad_dir;
    end
    if (sel) begin
      lineBuffer_220_value <= lineBuffer_219_value;
    end
    if (sel) begin
      lineBuffer_221_grad_dir <= lineBuffer_220_grad_dir;
    end
    if (sel) begin
      lineBuffer_221_value <= lineBuffer_220_value;
    end
    if (sel) begin
      lineBuffer_222_grad_dir <= lineBuffer_221_grad_dir;
    end
    if (sel) begin
      lineBuffer_222_value <= lineBuffer_221_value;
    end
    if (sel) begin
      lineBuffer_223_grad_dir <= lineBuffer_222_grad_dir;
    end
    if (sel) begin
      lineBuffer_223_value <= lineBuffer_222_value;
    end
    if (sel) begin
      lineBuffer_224_grad_dir <= lineBuffer_223_grad_dir;
    end
    if (sel) begin
      lineBuffer_224_value <= lineBuffer_223_value;
    end
    if (sel) begin
      lineBuffer_225_grad_dir <= lineBuffer_224_grad_dir;
    end
    if (sel) begin
      lineBuffer_225_value <= lineBuffer_224_value;
    end
    if (sel) begin
      lineBuffer_226_grad_dir <= lineBuffer_225_grad_dir;
    end
    if (sel) begin
      lineBuffer_226_value <= lineBuffer_225_value;
    end
    if (sel) begin
      lineBuffer_227_grad_dir <= lineBuffer_226_grad_dir;
    end
    if (sel) begin
      lineBuffer_227_value <= lineBuffer_226_value;
    end
    if (sel) begin
      lineBuffer_228_grad_dir <= lineBuffer_227_grad_dir;
    end
    if (sel) begin
      lineBuffer_228_value <= lineBuffer_227_value;
    end
    if (sel) begin
      lineBuffer_229_grad_dir <= lineBuffer_228_grad_dir;
    end
    if (sel) begin
      lineBuffer_229_value <= lineBuffer_228_value;
    end
    if (sel) begin
      lineBuffer_230_grad_dir <= lineBuffer_229_grad_dir;
    end
    if (sel) begin
      lineBuffer_230_value <= lineBuffer_229_value;
    end
    if (sel) begin
      lineBuffer_231_grad_dir <= lineBuffer_230_grad_dir;
    end
    if (sel) begin
      lineBuffer_231_value <= lineBuffer_230_value;
    end
    if (sel) begin
      lineBuffer_232_grad_dir <= lineBuffer_231_grad_dir;
    end
    if (sel) begin
      lineBuffer_232_value <= lineBuffer_231_value;
    end
    if (sel) begin
      lineBuffer_233_grad_dir <= lineBuffer_232_grad_dir;
    end
    if (sel) begin
      lineBuffer_233_value <= lineBuffer_232_value;
    end
    if (sel) begin
      lineBuffer_234_grad_dir <= lineBuffer_233_grad_dir;
    end
    if (sel) begin
      lineBuffer_234_value <= lineBuffer_233_value;
    end
    if (sel) begin
      lineBuffer_235_grad_dir <= lineBuffer_234_grad_dir;
    end
    if (sel) begin
      lineBuffer_235_value <= lineBuffer_234_value;
    end
    if (sel) begin
      lineBuffer_236_grad_dir <= lineBuffer_235_grad_dir;
    end
    if (sel) begin
      lineBuffer_236_value <= lineBuffer_235_value;
    end
    if (sel) begin
      lineBuffer_237_grad_dir <= lineBuffer_236_grad_dir;
    end
    if (sel) begin
      lineBuffer_237_value <= lineBuffer_236_value;
    end
    if (sel) begin
      lineBuffer_238_grad_dir <= lineBuffer_237_grad_dir;
    end
    if (sel) begin
      lineBuffer_238_value <= lineBuffer_237_value;
    end
    if (sel) begin
      lineBuffer_239_grad_dir <= lineBuffer_238_grad_dir;
    end
    if (sel) begin
      lineBuffer_239_value <= lineBuffer_238_value;
    end
    if (sel) begin
      lineBuffer_240_grad_dir <= lineBuffer_239_grad_dir;
    end
    if (sel) begin
      lineBuffer_240_value <= lineBuffer_239_value;
    end
    if (sel) begin
      lineBuffer_241_grad_dir <= lineBuffer_240_grad_dir;
    end
    if (sel) begin
      lineBuffer_241_value <= lineBuffer_240_value;
    end
    if (sel) begin
      lineBuffer_242_grad_dir <= lineBuffer_241_grad_dir;
    end
    if (sel) begin
      lineBuffer_242_value <= lineBuffer_241_value;
    end
    if (sel) begin
      lineBuffer_243_grad_dir <= lineBuffer_242_grad_dir;
    end
    if (sel) begin
      lineBuffer_243_value <= lineBuffer_242_value;
    end
    if (sel) begin
      lineBuffer_244_grad_dir <= lineBuffer_243_grad_dir;
    end
    if (sel) begin
      lineBuffer_244_value <= lineBuffer_243_value;
    end
    if (sel) begin
      lineBuffer_245_grad_dir <= lineBuffer_244_grad_dir;
    end
    if (sel) begin
      lineBuffer_245_value <= lineBuffer_244_value;
    end
    if (sel) begin
      lineBuffer_246_grad_dir <= lineBuffer_245_grad_dir;
    end
    if (sel) begin
      lineBuffer_246_value <= lineBuffer_245_value;
    end
    if (sel) begin
      lineBuffer_247_grad_dir <= lineBuffer_246_grad_dir;
    end
    if (sel) begin
      lineBuffer_247_value <= lineBuffer_246_value;
    end
    if (sel) begin
      lineBuffer_248_grad_dir <= lineBuffer_247_grad_dir;
    end
    if (sel) begin
      lineBuffer_248_value <= lineBuffer_247_value;
    end
    if (sel) begin
      lineBuffer_249_grad_dir <= lineBuffer_248_grad_dir;
    end
    if (sel) begin
      lineBuffer_249_value <= lineBuffer_248_value;
    end
    if (sel) begin
      lineBuffer_250_grad_dir <= lineBuffer_249_grad_dir;
    end
    if (sel) begin
      lineBuffer_250_value <= lineBuffer_249_value;
    end
    if (sel) begin
      lineBuffer_251_grad_dir <= lineBuffer_250_grad_dir;
    end
    if (sel) begin
      lineBuffer_251_value <= lineBuffer_250_value;
    end
    if (sel) begin
      lineBuffer_252_grad_dir <= lineBuffer_251_grad_dir;
    end
    if (sel) begin
      lineBuffer_252_value <= lineBuffer_251_value;
    end
    if (sel) begin
      lineBuffer_253_grad_dir <= lineBuffer_252_grad_dir;
    end
    if (sel) begin
      lineBuffer_253_value <= lineBuffer_252_value;
    end
    if (sel) begin
      lineBuffer_254_grad_dir <= lineBuffer_253_grad_dir;
    end
    if (sel) begin
      lineBuffer_254_value <= lineBuffer_253_value;
    end
    if (sel) begin
      lineBuffer_255_grad_dir <= lineBuffer_254_grad_dir;
    end
    if (sel) begin
      lineBuffer_255_value <= lineBuffer_254_value;
    end
    if (sel) begin
      lineBuffer_256_grad_dir <= lineBuffer_255_grad_dir;
    end
    if (sel) begin
      lineBuffer_256_value <= lineBuffer_255_value;
    end
    if (sel) begin
      lineBuffer_257_grad_dir <= lineBuffer_256_grad_dir;
    end
    if (sel) begin
      lineBuffer_257_value <= lineBuffer_256_value;
    end
    if (sel) begin
      lineBuffer_258_grad_dir <= lineBuffer_257_grad_dir;
    end
    if (sel) begin
      lineBuffer_258_value <= lineBuffer_257_value;
    end
    if (sel) begin
      lineBuffer_259_grad_dir <= lineBuffer_258_grad_dir;
    end
    if (sel) begin
      lineBuffer_259_value <= lineBuffer_258_value;
    end
    if (sel) begin
      lineBuffer_260_grad_dir <= lineBuffer_259_grad_dir;
    end
    if (sel) begin
      lineBuffer_260_value <= lineBuffer_259_value;
    end
    if (sel) begin
      lineBuffer_261_grad_dir <= lineBuffer_260_grad_dir;
    end
    if (sel) begin
      lineBuffer_261_value <= lineBuffer_260_value;
    end
    if (sel) begin
      lineBuffer_262_grad_dir <= lineBuffer_261_grad_dir;
    end
    if (sel) begin
      lineBuffer_262_value <= lineBuffer_261_value;
    end
    if (sel) begin
      lineBuffer_263_grad_dir <= lineBuffer_262_grad_dir;
    end
    if (sel) begin
      lineBuffer_263_value <= lineBuffer_262_value;
    end
    if (sel) begin
      lineBuffer_264_grad_dir <= lineBuffer_263_grad_dir;
    end
    if (sel) begin
      lineBuffer_264_value <= lineBuffer_263_value;
    end
    if (sel) begin
      lineBuffer_265_grad_dir <= lineBuffer_264_grad_dir;
    end
    if (sel) begin
      lineBuffer_265_value <= lineBuffer_264_value;
    end
    if (sel) begin
      lineBuffer_266_grad_dir <= lineBuffer_265_grad_dir;
    end
    if (sel) begin
      lineBuffer_266_value <= lineBuffer_265_value;
    end
    if (sel) begin
      lineBuffer_267_grad_dir <= lineBuffer_266_grad_dir;
    end
    if (sel) begin
      lineBuffer_267_value <= lineBuffer_266_value;
    end
    if (sel) begin
      lineBuffer_268_grad_dir <= lineBuffer_267_grad_dir;
    end
    if (sel) begin
      lineBuffer_268_value <= lineBuffer_267_value;
    end
    if (sel) begin
      lineBuffer_269_grad_dir <= lineBuffer_268_grad_dir;
    end
    if (sel) begin
      lineBuffer_269_value <= lineBuffer_268_value;
    end
    if (sel) begin
      lineBuffer_270_grad_dir <= lineBuffer_269_grad_dir;
    end
    if (sel) begin
      lineBuffer_270_value <= lineBuffer_269_value;
    end
    if (sel) begin
      lineBuffer_271_grad_dir <= lineBuffer_270_grad_dir;
    end
    if (sel) begin
      lineBuffer_271_value <= lineBuffer_270_value;
    end
    if (sel) begin
      lineBuffer_272_grad_dir <= lineBuffer_271_grad_dir;
    end
    if (sel) begin
      lineBuffer_272_value <= lineBuffer_271_value;
    end
    if (sel) begin
      lineBuffer_273_grad_dir <= lineBuffer_272_grad_dir;
    end
    if (sel) begin
      lineBuffer_273_value <= lineBuffer_272_value;
    end
    if (sel) begin
      lineBuffer_274_grad_dir <= lineBuffer_273_grad_dir;
    end
    if (sel) begin
      lineBuffer_274_value <= lineBuffer_273_value;
    end
    if (sel) begin
      lineBuffer_275_grad_dir <= lineBuffer_274_grad_dir;
    end
    if (sel) begin
      lineBuffer_275_value <= lineBuffer_274_value;
    end
    if (sel) begin
      lineBuffer_276_grad_dir <= lineBuffer_275_grad_dir;
    end
    if (sel) begin
      lineBuffer_276_value <= lineBuffer_275_value;
    end
    if (sel) begin
      lineBuffer_277_grad_dir <= lineBuffer_276_grad_dir;
    end
    if (sel) begin
      lineBuffer_277_value <= lineBuffer_276_value;
    end
    if (sel) begin
      lineBuffer_278_grad_dir <= lineBuffer_277_grad_dir;
    end
    if (sel) begin
      lineBuffer_278_value <= lineBuffer_277_value;
    end
    if (sel) begin
      lineBuffer_279_grad_dir <= lineBuffer_278_grad_dir;
    end
    if (sel) begin
      lineBuffer_279_value <= lineBuffer_278_value;
    end
    if (sel) begin
      lineBuffer_280_grad_dir <= lineBuffer_279_grad_dir;
    end
    if (sel) begin
      lineBuffer_280_value <= lineBuffer_279_value;
    end
    if (sel) begin
      lineBuffer_281_grad_dir <= lineBuffer_280_grad_dir;
    end
    if (sel) begin
      lineBuffer_281_value <= lineBuffer_280_value;
    end
    if (sel) begin
      lineBuffer_282_grad_dir <= lineBuffer_281_grad_dir;
    end
    if (sel) begin
      lineBuffer_282_value <= lineBuffer_281_value;
    end
    if (sel) begin
      lineBuffer_283_grad_dir <= lineBuffer_282_grad_dir;
    end
    if (sel) begin
      lineBuffer_283_value <= lineBuffer_282_value;
    end
    if (sel) begin
      lineBuffer_284_grad_dir <= lineBuffer_283_grad_dir;
    end
    if (sel) begin
      lineBuffer_284_value <= lineBuffer_283_value;
    end
    if (sel) begin
      lineBuffer_285_grad_dir <= lineBuffer_284_grad_dir;
    end
    if (sel) begin
      lineBuffer_285_value <= lineBuffer_284_value;
    end
    if (sel) begin
      lineBuffer_286_grad_dir <= lineBuffer_285_grad_dir;
    end
    if (sel) begin
      lineBuffer_286_value <= lineBuffer_285_value;
    end
    if (sel) begin
      lineBuffer_287_grad_dir <= lineBuffer_286_grad_dir;
    end
    if (sel) begin
      lineBuffer_287_value <= lineBuffer_286_value;
    end
    if (sel) begin
      lineBuffer_288_grad_dir <= lineBuffer_287_grad_dir;
    end
    if (sel) begin
      lineBuffer_288_value <= lineBuffer_287_value;
    end
    if (sel) begin
      lineBuffer_289_grad_dir <= lineBuffer_288_grad_dir;
    end
    if (sel) begin
      lineBuffer_289_value <= lineBuffer_288_value;
    end
    if (sel) begin
      lineBuffer_290_grad_dir <= lineBuffer_289_grad_dir;
    end
    if (sel) begin
      lineBuffer_290_value <= lineBuffer_289_value;
    end
    if (sel) begin
      lineBuffer_291_grad_dir <= lineBuffer_290_grad_dir;
    end
    if (sel) begin
      lineBuffer_291_value <= lineBuffer_290_value;
    end
    if (sel) begin
      lineBuffer_292_grad_dir <= lineBuffer_291_grad_dir;
    end
    if (sel) begin
      lineBuffer_292_value <= lineBuffer_291_value;
    end
    if (sel) begin
      lineBuffer_293_grad_dir <= lineBuffer_292_grad_dir;
    end
    if (sel) begin
      lineBuffer_293_value <= lineBuffer_292_value;
    end
    if (sel) begin
      lineBuffer_294_grad_dir <= lineBuffer_293_grad_dir;
    end
    if (sel) begin
      lineBuffer_294_value <= lineBuffer_293_value;
    end
    if (sel) begin
      lineBuffer_295_grad_dir <= lineBuffer_294_grad_dir;
    end
    if (sel) begin
      lineBuffer_295_value <= lineBuffer_294_value;
    end
    if (sel) begin
      lineBuffer_296_grad_dir <= lineBuffer_295_grad_dir;
    end
    if (sel) begin
      lineBuffer_296_value <= lineBuffer_295_value;
    end
    if (sel) begin
      lineBuffer_297_grad_dir <= lineBuffer_296_grad_dir;
    end
    if (sel) begin
      lineBuffer_297_value <= lineBuffer_296_value;
    end
    if (sel) begin
      lineBuffer_298_grad_dir <= lineBuffer_297_grad_dir;
    end
    if (sel) begin
      lineBuffer_298_value <= lineBuffer_297_value;
    end
    if (sel) begin
      lineBuffer_299_grad_dir <= lineBuffer_298_grad_dir;
    end
    if (sel) begin
      lineBuffer_299_value <= lineBuffer_298_value;
    end
    if (sel) begin
      lineBuffer_300_grad_dir <= lineBuffer_299_grad_dir;
    end
    if (sel) begin
      lineBuffer_300_value <= lineBuffer_299_value;
    end
    if (sel) begin
      lineBuffer_301_grad_dir <= lineBuffer_300_grad_dir;
    end
    if (sel) begin
      lineBuffer_301_value <= lineBuffer_300_value;
    end
    if (sel) begin
      lineBuffer_302_grad_dir <= lineBuffer_301_grad_dir;
    end
    if (sel) begin
      lineBuffer_302_value <= lineBuffer_301_value;
    end
    if (sel) begin
      lineBuffer_303_grad_dir <= lineBuffer_302_grad_dir;
    end
    if (sel) begin
      lineBuffer_303_value <= lineBuffer_302_value;
    end
    if (sel) begin
      lineBuffer_304_grad_dir <= lineBuffer_303_grad_dir;
    end
    if (sel) begin
      lineBuffer_304_value <= lineBuffer_303_value;
    end
    if (sel) begin
      lineBuffer_305_grad_dir <= lineBuffer_304_grad_dir;
    end
    if (sel) begin
      lineBuffer_305_value <= lineBuffer_304_value;
    end
    if (sel) begin
      lineBuffer_306_grad_dir <= lineBuffer_305_grad_dir;
    end
    if (sel) begin
      lineBuffer_306_value <= lineBuffer_305_value;
    end
    if (sel) begin
      lineBuffer_307_grad_dir <= lineBuffer_306_grad_dir;
    end
    if (sel) begin
      lineBuffer_307_value <= lineBuffer_306_value;
    end
    if (sel) begin
      lineBuffer_308_grad_dir <= lineBuffer_307_grad_dir;
    end
    if (sel) begin
      lineBuffer_308_value <= lineBuffer_307_value;
    end
    if (sel) begin
      lineBuffer_309_grad_dir <= lineBuffer_308_grad_dir;
    end
    if (sel) begin
      lineBuffer_309_value <= lineBuffer_308_value;
    end
    if (sel) begin
      lineBuffer_310_grad_dir <= lineBuffer_309_grad_dir;
    end
    if (sel) begin
      lineBuffer_310_value <= lineBuffer_309_value;
    end
    if (sel) begin
      lineBuffer_311_grad_dir <= lineBuffer_310_grad_dir;
    end
    if (sel) begin
      lineBuffer_311_value <= lineBuffer_310_value;
    end
    if (sel) begin
      lineBuffer_312_grad_dir <= lineBuffer_311_grad_dir;
    end
    if (sel) begin
      lineBuffer_312_value <= lineBuffer_311_value;
    end
    if (sel) begin
      lineBuffer_313_grad_dir <= lineBuffer_312_grad_dir;
    end
    if (sel) begin
      lineBuffer_313_value <= lineBuffer_312_value;
    end
    if (sel) begin
      lineBuffer_314_grad_dir <= lineBuffer_313_grad_dir;
    end
    if (sel) begin
      lineBuffer_314_value <= lineBuffer_313_value;
    end
    if (sel) begin
      lineBuffer_315_grad_dir <= lineBuffer_314_grad_dir;
    end
    if (sel) begin
      lineBuffer_315_value <= lineBuffer_314_value;
    end
    if (sel) begin
      lineBuffer_316_grad_dir <= lineBuffer_315_grad_dir;
    end
    if (sel) begin
      lineBuffer_316_value <= lineBuffer_315_value;
    end
    if (sel) begin
      lineBuffer_317_grad_dir <= lineBuffer_316_grad_dir;
    end
    if (sel) begin
      lineBuffer_317_value <= lineBuffer_316_value;
    end
    if (sel) begin
      lineBuffer_318_grad_dir <= lineBuffer_317_grad_dir;
    end
    if (sel) begin
      lineBuffer_318_value <= lineBuffer_317_value;
    end
    if (sel) begin
      lineBuffer_319_grad_dir <= lineBuffer_318_grad_dir;
    end
    if (sel) begin
      lineBuffer_319_value <= lineBuffer_318_value;
    end
    if (sel) begin
      lineBuffer_320_grad_dir <= lineBuffer_319_grad_dir;
    end
    if (sel) begin
      lineBuffer_320_value <= lineBuffer_319_value;
    end
    if (sel) begin
      lineBuffer_321_grad_dir <= lineBuffer_320_grad_dir;
    end
    if (sel) begin
      lineBuffer_321_value <= lineBuffer_320_value;
    end
    if (sel) begin
      lineBuffer_322_grad_dir <= lineBuffer_321_grad_dir;
    end
    if (sel) begin
      lineBuffer_322_value <= lineBuffer_321_value;
    end
    if (sel) begin
      lineBuffer_323_grad_dir <= lineBuffer_322_grad_dir;
    end
    if (sel) begin
      lineBuffer_323_value <= lineBuffer_322_value;
    end
    if (sel) begin
      lineBuffer_324_grad_dir <= lineBuffer_323_grad_dir;
    end
    if (sel) begin
      lineBuffer_324_value <= lineBuffer_323_value;
    end
    if (sel) begin
      lineBuffer_325_grad_dir <= lineBuffer_324_grad_dir;
    end
    if (sel) begin
      lineBuffer_325_value <= lineBuffer_324_value;
    end
    if (sel) begin
      lineBuffer_326_grad_dir <= lineBuffer_325_grad_dir;
    end
    if (sel) begin
      lineBuffer_326_value <= lineBuffer_325_value;
    end
    if (sel) begin
      lineBuffer_327_grad_dir <= lineBuffer_326_grad_dir;
    end
    if (sel) begin
      lineBuffer_327_value <= lineBuffer_326_value;
    end
    if (sel) begin
      lineBuffer_328_grad_dir <= lineBuffer_327_grad_dir;
    end
    if (sel) begin
      lineBuffer_328_value <= lineBuffer_327_value;
    end
    if (sel) begin
      lineBuffer_329_grad_dir <= lineBuffer_328_grad_dir;
    end
    if (sel) begin
      lineBuffer_329_value <= lineBuffer_328_value;
    end
    if (sel) begin
      lineBuffer_330_grad_dir <= lineBuffer_329_grad_dir;
    end
    if (sel) begin
      lineBuffer_330_value <= lineBuffer_329_value;
    end
    if (sel) begin
      lineBuffer_331_grad_dir <= lineBuffer_330_grad_dir;
    end
    if (sel) begin
      lineBuffer_331_value <= lineBuffer_330_value;
    end
    if (sel) begin
      lineBuffer_332_grad_dir <= lineBuffer_331_grad_dir;
    end
    if (sel) begin
      lineBuffer_332_value <= lineBuffer_331_value;
    end
    if (sel) begin
      lineBuffer_333_grad_dir <= lineBuffer_332_grad_dir;
    end
    if (sel) begin
      lineBuffer_333_value <= lineBuffer_332_value;
    end
    if (sel) begin
      lineBuffer_334_grad_dir <= lineBuffer_333_grad_dir;
    end
    if (sel) begin
      lineBuffer_334_value <= lineBuffer_333_value;
    end
    if (sel) begin
      lineBuffer_335_grad_dir <= lineBuffer_334_grad_dir;
    end
    if (sel) begin
      lineBuffer_335_value <= lineBuffer_334_value;
    end
    if (sel) begin
      lineBuffer_336_grad_dir <= lineBuffer_335_grad_dir;
    end
    if (sel) begin
      lineBuffer_336_value <= lineBuffer_335_value;
    end
    if (sel) begin
      lineBuffer_337_grad_dir <= lineBuffer_336_grad_dir;
    end
    if (sel) begin
      lineBuffer_337_value <= lineBuffer_336_value;
    end
    if (sel) begin
      lineBuffer_338_grad_dir <= lineBuffer_337_grad_dir;
    end
    if (sel) begin
      lineBuffer_338_value <= lineBuffer_337_value;
    end
    if (sel) begin
      lineBuffer_339_grad_dir <= lineBuffer_338_grad_dir;
    end
    if (sel) begin
      lineBuffer_339_value <= lineBuffer_338_value;
    end
    if (sel) begin
      lineBuffer_340_grad_dir <= lineBuffer_339_grad_dir;
    end
    if (sel) begin
      lineBuffer_340_value <= lineBuffer_339_value;
    end
    if (sel) begin
      lineBuffer_341_grad_dir <= lineBuffer_340_grad_dir;
    end
    if (sel) begin
      lineBuffer_341_value <= lineBuffer_340_value;
    end
    if (sel) begin
      lineBuffer_342_grad_dir <= lineBuffer_341_grad_dir;
    end
    if (sel) begin
      lineBuffer_342_value <= lineBuffer_341_value;
    end
    if (sel) begin
      lineBuffer_343_grad_dir <= lineBuffer_342_grad_dir;
    end
    if (sel) begin
      lineBuffer_343_value <= lineBuffer_342_value;
    end
    if (sel) begin
      lineBuffer_344_grad_dir <= lineBuffer_343_grad_dir;
    end
    if (sel) begin
      lineBuffer_344_value <= lineBuffer_343_value;
    end
    if (sel) begin
      lineBuffer_345_grad_dir <= lineBuffer_344_grad_dir;
    end
    if (sel) begin
      lineBuffer_345_value <= lineBuffer_344_value;
    end
    if (sel) begin
      lineBuffer_346_grad_dir <= lineBuffer_345_grad_dir;
    end
    if (sel) begin
      lineBuffer_346_value <= lineBuffer_345_value;
    end
    if (sel) begin
      lineBuffer_347_grad_dir <= lineBuffer_346_grad_dir;
    end
    if (sel) begin
      lineBuffer_347_value <= lineBuffer_346_value;
    end
    if (sel) begin
      lineBuffer_348_grad_dir <= lineBuffer_347_grad_dir;
    end
    if (sel) begin
      lineBuffer_348_value <= lineBuffer_347_value;
    end
    if (sel) begin
      lineBuffer_349_grad_dir <= lineBuffer_348_grad_dir;
    end
    if (sel) begin
      lineBuffer_349_value <= lineBuffer_348_value;
    end
    if (sel) begin
      lineBuffer_350_grad_dir <= lineBuffer_349_grad_dir;
    end
    if (sel) begin
      lineBuffer_350_value <= lineBuffer_349_value;
    end
    if (sel) begin
      lineBuffer_351_grad_dir <= lineBuffer_350_grad_dir;
    end
    if (sel) begin
      lineBuffer_351_value <= lineBuffer_350_value;
    end
    if (sel) begin
      lineBuffer_352_grad_dir <= lineBuffer_351_grad_dir;
    end
    if (sel) begin
      lineBuffer_352_value <= lineBuffer_351_value;
    end
    if (sel) begin
      lineBuffer_353_grad_dir <= lineBuffer_352_grad_dir;
    end
    if (sel) begin
      lineBuffer_353_value <= lineBuffer_352_value;
    end
    if (sel) begin
      lineBuffer_354_grad_dir <= lineBuffer_353_grad_dir;
    end
    if (sel) begin
      lineBuffer_354_value <= lineBuffer_353_value;
    end
    if (sel) begin
      lineBuffer_355_grad_dir <= lineBuffer_354_grad_dir;
    end
    if (sel) begin
      lineBuffer_355_value <= lineBuffer_354_value;
    end
    if (sel) begin
      lineBuffer_356_grad_dir <= lineBuffer_355_grad_dir;
    end
    if (sel) begin
      lineBuffer_356_value <= lineBuffer_355_value;
    end
    if (sel) begin
      lineBuffer_357_grad_dir <= lineBuffer_356_grad_dir;
    end
    if (sel) begin
      lineBuffer_357_value <= lineBuffer_356_value;
    end
    if (sel) begin
      lineBuffer_358_grad_dir <= lineBuffer_357_grad_dir;
    end
    if (sel) begin
      lineBuffer_358_value <= lineBuffer_357_value;
    end
    if (sel) begin
      lineBuffer_359_grad_dir <= lineBuffer_358_grad_dir;
    end
    if (sel) begin
      lineBuffer_359_value <= lineBuffer_358_value;
    end
    if (sel) begin
      lineBuffer_360_grad_dir <= lineBuffer_359_grad_dir;
    end
    if (sel) begin
      lineBuffer_360_value <= lineBuffer_359_value;
    end
    if (sel) begin
      lineBuffer_361_grad_dir <= lineBuffer_360_grad_dir;
    end
    if (sel) begin
      lineBuffer_361_value <= lineBuffer_360_value;
    end
    if (sel) begin
      lineBuffer_362_grad_dir <= lineBuffer_361_grad_dir;
    end
    if (sel) begin
      lineBuffer_362_value <= lineBuffer_361_value;
    end
    if (sel) begin
      lineBuffer_363_grad_dir <= lineBuffer_362_grad_dir;
    end
    if (sel) begin
      lineBuffer_363_value <= lineBuffer_362_value;
    end
    if (sel) begin
      lineBuffer_364_grad_dir <= lineBuffer_363_grad_dir;
    end
    if (sel) begin
      lineBuffer_364_value <= lineBuffer_363_value;
    end
    if (sel) begin
      lineBuffer_365_grad_dir <= lineBuffer_364_grad_dir;
    end
    if (sel) begin
      lineBuffer_365_value <= lineBuffer_364_value;
    end
    if (sel) begin
      lineBuffer_366_grad_dir <= lineBuffer_365_grad_dir;
    end
    if (sel) begin
      lineBuffer_366_value <= lineBuffer_365_value;
    end
    if (sel) begin
      lineBuffer_367_grad_dir <= lineBuffer_366_grad_dir;
    end
    if (sel) begin
      lineBuffer_367_value <= lineBuffer_366_value;
    end
    if (sel) begin
      lineBuffer_368_grad_dir <= lineBuffer_367_grad_dir;
    end
    if (sel) begin
      lineBuffer_368_value <= lineBuffer_367_value;
    end
    if (sel) begin
      lineBuffer_369_grad_dir <= lineBuffer_368_grad_dir;
    end
    if (sel) begin
      lineBuffer_369_value <= lineBuffer_368_value;
    end
    if (sel) begin
      lineBuffer_370_grad_dir <= lineBuffer_369_grad_dir;
    end
    if (sel) begin
      lineBuffer_370_value <= lineBuffer_369_value;
    end
    if (sel) begin
      lineBuffer_371_grad_dir <= lineBuffer_370_grad_dir;
    end
    if (sel) begin
      lineBuffer_371_value <= lineBuffer_370_value;
    end
    if (sel) begin
      lineBuffer_372_grad_dir <= lineBuffer_371_grad_dir;
    end
    if (sel) begin
      lineBuffer_372_value <= lineBuffer_371_value;
    end
    if (sel) begin
      lineBuffer_373_grad_dir <= lineBuffer_372_grad_dir;
    end
    if (sel) begin
      lineBuffer_373_value <= lineBuffer_372_value;
    end
    if (sel) begin
      lineBuffer_374_grad_dir <= lineBuffer_373_grad_dir;
    end
    if (sel) begin
      lineBuffer_374_value <= lineBuffer_373_value;
    end
    if (sel) begin
      lineBuffer_375_grad_dir <= lineBuffer_374_grad_dir;
    end
    if (sel) begin
      lineBuffer_375_value <= lineBuffer_374_value;
    end
    if (sel) begin
      lineBuffer_376_grad_dir <= lineBuffer_375_grad_dir;
    end
    if (sel) begin
      lineBuffer_376_value <= lineBuffer_375_value;
    end
    if (sel) begin
      lineBuffer_377_grad_dir <= lineBuffer_376_grad_dir;
    end
    if (sel) begin
      lineBuffer_377_value <= lineBuffer_376_value;
    end
    if (sel) begin
      lineBuffer_378_grad_dir <= lineBuffer_377_grad_dir;
    end
    if (sel) begin
      lineBuffer_378_value <= lineBuffer_377_value;
    end
    if (sel) begin
      lineBuffer_379_grad_dir <= lineBuffer_378_grad_dir;
    end
    if (sel) begin
      lineBuffer_379_value <= lineBuffer_378_value;
    end
    if (sel) begin
      lineBuffer_380_grad_dir <= lineBuffer_379_grad_dir;
    end
    if (sel) begin
      lineBuffer_380_value <= lineBuffer_379_value;
    end
    if (sel) begin
      lineBuffer_381_grad_dir <= lineBuffer_380_grad_dir;
    end
    if (sel) begin
      lineBuffer_381_value <= lineBuffer_380_value;
    end
    if (sel) begin
      lineBuffer_382_grad_dir <= lineBuffer_381_grad_dir;
    end
    if (sel) begin
      lineBuffer_382_value <= lineBuffer_381_value;
    end
    if (sel) begin
      lineBuffer_383_grad_dir <= lineBuffer_382_grad_dir;
    end
    if (sel) begin
      lineBuffer_383_value <= lineBuffer_382_value;
    end
    if (sel) begin
      lineBuffer_384_grad_dir <= lineBuffer_383_grad_dir;
    end
    if (sel) begin
      lineBuffer_384_value <= lineBuffer_383_value;
    end
    if (sel) begin
      lineBuffer_385_grad_dir <= lineBuffer_384_grad_dir;
    end
    if (sel) begin
      lineBuffer_385_value <= lineBuffer_384_value;
    end
    if (sel) begin
      lineBuffer_386_grad_dir <= lineBuffer_385_grad_dir;
    end
    if (sel) begin
      lineBuffer_386_value <= lineBuffer_385_value;
    end
    if (sel) begin
      lineBuffer_387_grad_dir <= lineBuffer_386_grad_dir;
    end
    if (sel) begin
      lineBuffer_387_value <= lineBuffer_386_value;
    end
    if (sel) begin
      lineBuffer_388_grad_dir <= lineBuffer_387_grad_dir;
    end
    if (sel) begin
      lineBuffer_388_value <= lineBuffer_387_value;
    end
    if (sel) begin
      lineBuffer_389_grad_dir <= lineBuffer_388_grad_dir;
    end
    if (sel) begin
      lineBuffer_389_value <= lineBuffer_388_value;
    end
    if (sel) begin
      lineBuffer_390_grad_dir <= lineBuffer_389_grad_dir;
    end
    if (sel) begin
      lineBuffer_390_value <= lineBuffer_389_value;
    end
    if (sel) begin
      lineBuffer_391_grad_dir <= lineBuffer_390_grad_dir;
    end
    if (sel) begin
      lineBuffer_391_value <= lineBuffer_390_value;
    end
    if (sel) begin
      lineBuffer_392_grad_dir <= lineBuffer_391_grad_dir;
    end
    if (sel) begin
      lineBuffer_392_value <= lineBuffer_391_value;
    end
    if (sel) begin
      lineBuffer_393_grad_dir <= lineBuffer_392_grad_dir;
    end
    if (sel) begin
      lineBuffer_393_value <= lineBuffer_392_value;
    end
    if (sel) begin
      lineBuffer_394_grad_dir <= lineBuffer_393_grad_dir;
    end
    if (sel) begin
      lineBuffer_394_value <= lineBuffer_393_value;
    end
    if (sel) begin
      lineBuffer_395_grad_dir <= lineBuffer_394_grad_dir;
    end
    if (sel) begin
      lineBuffer_395_value <= lineBuffer_394_value;
    end
    if (sel) begin
      lineBuffer_396_grad_dir <= lineBuffer_395_grad_dir;
    end
    if (sel) begin
      lineBuffer_396_value <= lineBuffer_395_value;
    end
    if (sel) begin
      lineBuffer_397_grad_dir <= lineBuffer_396_grad_dir;
    end
    if (sel) begin
      lineBuffer_397_value <= lineBuffer_396_value;
    end
    if (sel) begin
      lineBuffer_398_grad_dir <= lineBuffer_397_grad_dir;
    end
    if (sel) begin
      lineBuffer_398_value <= lineBuffer_397_value;
    end
    if (sel) begin
      lineBuffer_399_grad_dir <= lineBuffer_398_grad_dir;
    end
    if (sel) begin
      lineBuffer_399_value <= lineBuffer_398_value;
    end
    if (sel) begin
      lineBuffer_400_grad_dir <= lineBuffer_399_grad_dir;
    end
    if (sel) begin
      lineBuffer_400_value <= lineBuffer_399_value;
    end
    if (sel) begin
      lineBuffer_401_grad_dir <= lineBuffer_400_grad_dir;
    end
    if (sel) begin
      lineBuffer_401_value <= lineBuffer_400_value;
    end
    if (sel) begin
      lineBuffer_402_grad_dir <= lineBuffer_401_grad_dir;
    end
    if (sel) begin
      lineBuffer_402_value <= lineBuffer_401_value;
    end
    if (sel) begin
      lineBuffer_403_grad_dir <= lineBuffer_402_grad_dir;
    end
    if (sel) begin
      lineBuffer_403_value <= lineBuffer_402_value;
    end
    if (sel) begin
      lineBuffer_404_grad_dir <= lineBuffer_403_grad_dir;
    end
    if (sel) begin
      lineBuffer_404_value <= lineBuffer_403_value;
    end
    if (sel) begin
      lineBuffer_405_grad_dir <= lineBuffer_404_grad_dir;
    end
    if (sel) begin
      lineBuffer_405_value <= lineBuffer_404_value;
    end
    if (sel) begin
      lineBuffer_406_grad_dir <= lineBuffer_405_grad_dir;
    end
    if (sel) begin
      lineBuffer_406_value <= lineBuffer_405_value;
    end
    if (sel) begin
      lineBuffer_407_grad_dir <= lineBuffer_406_grad_dir;
    end
    if (sel) begin
      lineBuffer_407_value <= lineBuffer_406_value;
    end
    if (sel) begin
      lineBuffer_408_grad_dir <= lineBuffer_407_grad_dir;
    end
    if (sel) begin
      lineBuffer_408_value <= lineBuffer_407_value;
    end
    if (sel) begin
      lineBuffer_409_grad_dir <= lineBuffer_408_grad_dir;
    end
    if (sel) begin
      lineBuffer_409_value <= lineBuffer_408_value;
    end
    if (sel) begin
      lineBuffer_410_grad_dir <= lineBuffer_409_grad_dir;
    end
    if (sel) begin
      lineBuffer_410_value <= lineBuffer_409_value;
    end
    if (sel) begin
      lineBuffer_411_grad_dir <= lineBuffer_410_grad_dir;
    end
    if (sel) begin
      lineBuffer_411_value <= lineBuffer_410_value;
    end
    if (sel) begin
      lineBuffer_412_grad_dir <= lineBuffer_411_grad_dir;
    end
    if (sel) begin
      lineBuffer_412_value <= lineBuffer_411_value;
    end
    if (sel) begin
      lineBuffer_413_grad_dir <= lineBuffer_412_grad_dir;
    end
    if (sel) begin
      lineBuffer_413_value <= lineBuffer_412_value;
    end
    if (sel) begin
      lineBuffer_414_grad_dir <= lineBuffer_413_grad_dir;
    end
    if (sel) begin
      lineBuffer_414_value <= lineBuffer_413_value;
    end
    if (sel) begin
      lineBuffer_415_grad_dir <= lineBuffer_414_grad_dir;
    end
    if (sel) begin
      lineBuffer_415_value <= lineBuffer_414_value;
    end
    if (sel) begin
      lineBuffer_416_grad_dir <= lineBuffer_415_grad_dir;
    end
    if (sel) begin
      lineBuffer_416_value <= lineBuffer_415_value;
    end
    if (sel) begin
      lineBuffer_417_grad_dir <= lineBuffer_416_grad_dir;
    end
    if (sel) begin
      lineBuffer_417_value <= lineBuffer_416_value;
    end
    if (sel) begin
      lineBuffer_418_grad_dir <= lineBuffer_417_grad_dir;
    end
    if (sel) begin
      lineBuffer_418_value <= lineBuffer_417_value;
    end
    if (sel) begin
      lineBuffer_419_grad_dir <= lineBuffer_418_grad_dir;
    end
    if (sel) begin
      lineBuffer_419_value <= lineBuffer_418_value;
    end
    if (sel) begin
      lineBuffer_420_grad_dir <= lineBuffer_419_grad_dir;
    end
    if (sel) begin
      lineBuffer_420_value <= lineBuffer_419_value;
    end
    if (sel) begin
      lineBuffer_421_grad_dir <= lineBuffer_420_grad_dir;
    end
    if (sel) begin
      lineBuffer_421_value <= lineBuffer_420_value;
    end
    if (sel) begin
      lineBuffer_422_grad_dir <= lineBuffer_421_grad_dir;
    end
    if (sel) begin
      lineBuffer_422_value <= lineBuffer_421_value;
    end
    if (sel) begin
      lineBuffer_423_grad_dir <= lineBuffer_422_grad_dir;
    end
    if (sel) begin
      lineBuffer_423_value <= lineBuffer_422_value;
    end
    if (sel) begin
      lineBuffer_424_grad_dir <= lineBuffer_423_grad_dir;
    end
    if (sel) begin
      lineBuffer_424_value <= lineBuffer_423_value;
    end
    if (sel) begin
      lineBuffer_425_grad_dir <= lineBuffer_424_grad_dir;
    end
    if (sel) begin
      lineBuffer_425_value <= lineBuffer_424_value;
    end
    if (sel) begin
      lineBuffer_426_grad_dir <= lineBuffer_425_grad_dir;
    end
    if (sel) begin
      lineBuffer_426_value <= lineBuffer_425_value;
    end
    if (sel) begin
      lineBuffer_427_grad_dir <= lineBuffer_426_grad_dir;
    end
    if (sel) begin
      lineBuffer_427_value <= lineBuffer_426_value;
    end
    if (sel) begin
      lineBuffer_428_grad_dir <= lineBuffer_427_grad_dir;
    end
    if (sel) begin
      lineBuffer_428_value <= lineBuffer_427_value;
    end
    if (sel) begin
      lineBuffer_429_grad_dir <= lineBuffer_428_grad_dir;
    end
    if (sel) begin
      lineBuffer_429_value <= lineBuffer_428_value;
    end
    if (sel) begin
      lineBuffer_430_grad_dir <= lineBuffer_429_grad_dir;
    end
    if (sel) begin
      lineBuffer_430_value <= lineBuffer_429_value;
    end
    if (sel) begin
      lineBuffer_431_grad_dir <= lineBuffer_430_grad_dir;
    end
    if (sel) begin
      lineBuffer_431_value <= lineBuffer_430_value;
    end
    if (sel) begin
      lineBuffer_432_grad_dir <= lineBuffer_431_grad_dir;
    end
    if (sel) begin
      lineBuffer_432_value <= lineBuffer_431_value;
    end
    if (sel) begin
      lineBuffer_433_grad_dir <= lineBuffer_432_grad_dir;
    end
    if (sel) begin
      lineBuffer_433_value <= lineBuffer_432_value;
    end
    if (sel) begin
      lineBuffer_434_grad_dir <= lineBuffer_433_grad_dir;
    end
    if (sel) begin
      lineBuffer_434_value <= lineBuffer_433_value;
    end
    if (sel) begin
      lineBuffer_435_grad_dir <= lineBuffer_434_grad_dir;
    end
    if (sel) begin
      lineBuffer_435_value <= lineBuffer_434_value;
    end
    if (sel) begin
      lineBuffer_436_grad_dir <= lineBuffer_435_grad_dir;
    end
    if (sel) begin
      lineBuffer_436_value <= lineBuffer_435_value;
    end
    if (sel) begin
      lineBuffer_437_grad_dir <= lineBuffer_436_grad_dir;
    end
    if (sel) begin
      lineBuffer_437_value <= lineBuffer_436_value;
    end
    if (sel) begin
      lineBuffer_438_grad_dir <= lineBuffer_437_grad_dir;
    end
    if (sel) begin
      lineBuffer_438_value <= lineBuffer_437_value;
    end
    if (sel) begin
      lineBuffer_439_grad_dir <= lineBuffer_438_grad_dir;
    end
    if (sel) begin
      lineBuffer_439_value <= lineBuffer_438_value;
    end
    if (sel) begin
      lineBuffer_440_grad_dir <= lineBuffer_439_grad_dir;
    end
    if (sel) begin
      lineBuffer_440_value <= lineBuffer_439_value;
    end
    if (sel) begin
      lineBuffer_441_grad_dir <= lineBuffer_440_grad_dir;
    end
    if (sel) begin
      lineBuffer_441_value <= lineBuffer_440_value;
    end
    if (sel) begin
      lineBuffer_442_grad_dir <= lineBuffer_441_grad_dir;
    end
    if (sel) begin
      lineBuffer_442_value <= lineBuffer_441_value;
    end
    if (sel) begin
      lineBuffer_443_grad_dir <= lineBuffer_442_grad_dir;
    end
    if (sel) begin
      lineBuffer_443_value <= lineBuffer_442_value;
    end
    if (sel) begin
      lineBuffer_444_grad_dir <= lineBuffer_443_grad_dir;
    end
    if (sel) begin
      lineBuffer_444_value <= lineBuffer_443_value;
    end
    if (sel) begin
      lineBuffer_445_grad_dir <= lineBuffer_444_grad_dir;
    end
    if (sel) begin
      lineBuffer_445_value <= lineBuffer_444_value;
    end
    if (sel) begin
      lineBuffer_446_grad_dir <= lineBuffer_445_grad_dir;
    end
    if (sel) begin
      lineBuffer_446_value <= lineBuffer_445_value;
    end
    if (sel) begin
      lineBuffer_447_grad_dir <= lineBuffer_446_grad_dir;
    end
    if (sel) begin
      lineBuffer_447_value <= lineBuffer_446_value;
    end
    if (sel) begin
      lineBuffer_448_grad_dir <= lineBuffer_447_grad_dir;
    end
    if (sel) begin
      lineBuffer_448_value <= lineBuffer_447_value;
    end
    if (sel) begin
      lineBuffer_449_grad_dir <= lineBuffer_448_grad_dir;
    end
    if (sel) begin
      lineBuffer_449_value <= lineBuffer_448_value;
    end
    if (sel) begin
      lineBuffer_450_grad_dir <= lineBuffer_449_grad_dir;
    end
    if (sel) begin
      lineBuffer_450_value <= lineBuffer_449_value;
    end
    if (sel) begin
      lineBuffer_451_grad_dir <= lineBuffer_450_grad_dir;
    end
    if (sel) begin
      lineBuffer_451_value <= lineBuffer_450_value;
    end
    if (sel) begin
      lineBuffer_452_grad_dir <= lineBuffer_451_grad_dir;
    end
    if (sel) begin
      lineBuffer_452_value <= lineBuffer_451_value;
    end
    if (sel) begin
      lineBuffer_453_grad_dir <= lineBuffer_452_grad_dir;
    end
    if (sel) begin
      lineBuffer_453_value <= lineBuffer_452_value;
    end
    if (sel) begin
      lineBuffer_454_grad_dir <= lineBuffer_453_grad_dir;
    end
    if (sel) begin
      lineBuffer_454_value <= lineBuffer_453_value;
    end
    if (sel) begin
      lineBuffer_455_grad_dir <= lineBuffer_454_grad_dir;
    end
    if (sel) begin
      lineBuffer_455_value <= lineBuffer_454_value;
    end
    if (sel) begin
      lineBuffer_456_grad_dir <= lineBuffer_455_grad_dir;
    end
    if (sel) begin
      lineBuffer_456_value <= lineBuffer_455_value;
    end
    if (sel) begin
      lineBuffer_457_grad_dir <= lineBuffer_456_grad_dir;
    end
    if (sel) begin
      lineBuffer_457_value <= lineBuffer_456_value;
    end
    if (sel) begin
      lineBuffer_458_grad_dir <= lineBuffer_457_grad_dir;
    end
    if (sel) begin
      lineBuffer_458_value <= lineBuffer_457_value;
    end
    if (sel) begin
      lineBuffer_459_grad_dir <= lineBuffer_458_grad_dir;
    end
    if (sel) begin
      lineBuffer_459_value <= lineBuffer_458_value;
    end
    if (sel) begin
      lineBuffer_460_grad_dir <= lineBuffer_459_grad_dir;
    end
    if (sel) begin
      lineBuffer_460_value <= lineBuffer_459_value;
    end
    if (sel) begin
      lineBuffer_461_grad_dir <= lineBuffer_460_grad_dir;
    end
    if (sel) begin
      lineBuffer_461_value <= lineBuffer_460_value;
    end
    if (sel) begin
      lineBuffer_462_grad_dir <= lineBuffer_461_grad_dir;
    end
    if (sel) begin
      lineBuffer_462_value <= lineBuffer_461_value;
    end
    if (sel) begin
      lineBuffer_463_grad_dir <= lineBuffer_462_grad_dir;
    end
    if (sel) begin
      lineBuffer_463_value <= lineBuffer_462_value;
    end
    if (sel) begin
      lineBuffer_464_grad_dir <= lineBuffer_463_grad_dir;
    end
    if (sel) begin
      lineBuffer_464_value <= lineBuffer_463_value;
    end
    if (sel) begin
      lineBuffer_465_grad_dir <= lineBuffer_464_grad_dir;
    end
    if (sel) begin
      lineBuffer_465_value <= lineBuffer_464_value;
    end
    if (sel) begin
      lineBuffer_466_grad_dir <= lineBuffer_465_grad_dir;
    end
    if (sel) begin
      lineBuffer_466_value <= lineBuffer_465_value;
    end
    if (sel) begin
      lineBuffer_467_grad_dir <= lineBuffer_466_grad_dir;
    end
    if (sel) begin
      lineBuffer_467_value <= lineBuffer_466_value;
    end
    if (sel) begin
      lineBuffer_468_grad_dir <= lineBuffer_467_grad_dir;
    end
    if (sel) begin
      lineBuffer_468_value <= lineBuffer_467_value;
    end
    if (sel) begin
      lineBuffer_469_grad_dir <= lineBuffer_468_grad_dir;
    end
    if (sel) begin
      lineBuffer_469_value <= lineBuffer_468_value;
    end
    if (sel) begin
      lineBuffer_470_grad_dir <= lineBuffer_469_grad_dir;
    end
    if (sel) begin
      lineBuffer_470_value <= lineBuffer_469_value;
    end
    if (sel) begin
      lineBuffer_471_grad_dir <= lineBuffer_470_grad_dir;
    end
    if (sel) begin
      lineBuffer_471_value <= lineBuffer_470_value;
    end
    if (sel) begin
      lineBuffer_472_grad_dir <= lineBuffer_471_grad_dir;
    end
    if (sel) begin
      lineBuffer_472_value <= lineBuffer_471_value;
    end
    if (sel) begin
      lineBuffer_473_grad_dir <= lineBuffer_472_grad_dir;
    end
    if (sel) begin
      lineBuffer_473_value <= lineBuffer_472_value;
    end
    if (sel) begin
      lineBuffer_474_grad_dir <= lineBuffer_473_grad_dir;
    end
    if (sel) begin
      lineBuffer_474_value <= lineBuffer_473_value;
    end
    if (sel) begin
      lineBuffer_475_grad_dir <= lineBuffer_474_grad_dir;
    end
    if (sel) begin
      lineBuffer_475_value <= lineBuffer_474_value;
    end
    if (sel) begin
      lineBuffer_476_grad_dir <= lineBuffer_475_grad_dir;
    end
    if (sel) begin
      lineBuffer_476_value <= lineBuffer_475_value;
    end
    if (sel) begin
      lineBuffer_477_grad_dir <= lineBuffer_476_grad_dir;
    end
    if (sel) begin
      lineBuffer_477_value <= lineBuffer_476_value;
    end
    if (sel) begin
      lineBuffer_478_grad_dir <= lineBuffer_477_grad_dir;
    end
    if (sel) begin
      lineBuffer_478_value <= lineBuffer_477_value;
    end
    if (sel) begin
      lineBuffer_479_grad_dir <= lineBuffer_478_grad_dir;
    end
    if (sel) begin
      lineBuffer_479_value <= lineBuffer_478_value;
    end
    if (sel) begin
      lineBuffer_480_grad_dir <= lineBuffer_479_grad_dir;
    end
    if (sel) begin
      lineBuffer_480_value <= lineBuffer_479_value;
    end
    if (sel) begin
      lineBuffer_481_grad_dir <= lineBuffer_480_grad_dir;
    end
    if (sel) begin
      lineBuffer_481_value <= lineBuffer_480_value;
    end
    if (sel) begin
      lineBuffer_482_grad_dir <= lineBuffer_481_grad_dir;
    end
    if (sel) begin
      lineBuffer_482_value <= lineBuffer_481_value;
    end
    if (sel) begin
      lineBuffer_483_grad_dir <= lineBuffer_482_grad_dir;
    end
    if (sel) begin
      lineBuffer_483_value <= lineBuffer_482_value;
    end
    if (sel) begin
      lineBuffer_484_grad_dir <= lineBuffer_483_grad_dir;
    end
    if (sel) begin
      lineBuffer_484_value <= lineBuffer_483_value;
    end
    if (sel) begin
      lineBuffer_485_grad_dir <= lineBuffer_484_grad_dir;
    end
    if (sel) begin
      lineBuffer_485_value <= lineBuffer_484_value;
    end
    if (sel) begin
      lineBuffer_486_grad_dir <= lineBuffer_485_grad_dir;
    end
    if (sel) begin
      lineBuffer_486_value <= lineBuffer_485_value;
    end
    if (sel) begin
      lineBuffer_487_grad_dir <= lineBuffer_486_grad_dir;
    end
    if (sel) begin
      lineBuffer_487_value <= lineBuffer_486_value;
    end
    if (sel) begin
      lineBuffer_488_grad_dir <= lineBuffer_487_grad_dir;
    end
    if (sel) begin
      lineBuffer_488_value <= lineBuffer_487_value;
    end
    if (sel) begin
      lineBuffer_489_grad_dir <= lineBuffer_488_grad_dir;
    end
    if (sel) begin
      lineBuffer_489_value <= lineBuffer_488_value;
    end
    if (sel) begin
      lineBuffer_490_grad_dir <= lineBuffer_489_grad_dir;
    end
    if (sel) begin
      lineBuffer_490_value <= lineBuffer_489_value;
    end
    if (sel) begin
      lineBuffer_491_grad_dir <= lineBuffer_490_grad_dir;
    end
    if (sel) begin
      lineBuffer_491_value <= lineBuffer_490_value;
    end
    if (sel) begin
      lineBuffer_492_grad_dir <= lineBuffer_491_grad_dir;
    end
    if (sel) begin
      lineBuffer_492_value <= lineBuffer_491_value;
    end
    if (sel) begin
      lineBuffer_493_grad_dir <= lineBuffer_492_grad_dir;
    end
    if (sel) begin
      lineBuffer_493_value <= lineBuffer_492_value;
    end
    if (sel) begin
      lineBuffer_494_grad_dir <= lineBuffer_493_grad_dir;
    end
    if (sel) begin
      lineBuffer_494_value <= lineBuffer_493_value;
    end
    if (sel) begin
      lineBuffer_495_grad_dir <= lineBuffer_494_grad_dir;
    end
    if (sel) begin
      lineBuffer_495_value <= lineBuffer_494_value;
    end
    if (sel) begin
      lineBuffer_496_grad_dir <= lineBuffer_495_grad_dir;
    end
    if (sel) begin
      lineBuffer_496_value <= lineBuffer_495_value;
    end
    if (sel) begin
      lineBuffer_497_grad_dir <= lineBuffer_496_grad_dir;
    end
    if (sel) begin
      lineBuffer_497_value <= lineBuffer_496_value;
    end
    if (sel) begin
      lineBuffer_498_grad_dir <= lineBuffer_497_grad_dir;
    end
    if (sel) begin
      lineBuffer_498_value <= lineBuffer_497_value;
    end
    if (sel) begin
      lineBuffer_499_grad_dir <= lineBuffer_498_grad_dir;
    end
    if (sel) begin
      lineBuffer_499_value <= lineBuffer_498_value;
    end
    if (sel) begin
      lineBuffer_500_grad_dir <= lineBuffer_499_grad_dir;
    end
    if (sel) begin
      lineBuffer_500_value <= lineBuffer_499_value;
    end
    if (sel) begin
      lineBuffer_501_grad_dir <= lineBuffer_500_grad_dir;
    end
    if (sel) begin
      lineBuffer_501_value <= lineBuffer_500_value;
    end
    if (sel) begin
      lineBuffer_502_grad_dir <= lineBuffer_501_grad_dir;
    end
    if (sel) begin
      lineBuffer_502_value <= lineBuffer_501_value;
    end
    if (sel) begin
      lineBuffer_503_grad_dir <= lineBuffer_502_grad_dir;
    end
    if (sel) begin
      lineBuffer_503_value <= lineBuffer_502_value;
    end
    if (sel) begin
      lineBuffer_504_grad_dir <= lineBuffer_503_grad_dir;
    end
    if (sel) begin
      lineBuffer_504_value <= lineBuffer_503_value;
    end
    if (sel) begin
      lineBuffer_505_grad_dir <= lineBuffer_504_grad_dir;
    end
    if (sel) begin
      lineBuffer_505_value <= lineBuffer_504_value;
    end
    if (sel) begin
      lineBuffer_506_grad_dir <= lineBuffer_505_grad_dir;
    end
    if (sel) begin
      lineBuffer_506_value <= lineBuffer_505_value;
    end
    if (sel) begin
      lineBuffer_507_grad_dir <= lineBuffer_506_grad_dir;
    end
    if (sel) begin
      lineBuffer_507_value <= lineBuffer_506_value;
    end
    if (sel) begin
      lineBuffer_508_grad_dir <= lineBuffer_507_grad_dir;
    end
    if (sel) begin
      lineBuffer_508_value <= lineBuffer_507_value;
    end
    if (sel) begin
      lineBuffer_509_grad_dir <= lineBuffer_508_grad_dir;
    end
    if (sel) begin
      lineBuffer_509_value <= lineBuffer_508_value;
    end
    if (sel) begin
      lineBuffer_510_grad_dir <= lineBuffer_509_grad_dir;
    end
    if (sel) begin
      lineBuffer_510_value <= lineBuffer_509_value;
    end
    if (sel) begin
      lineBuffer_511_grad_dir <= lineBuffer_510_grad_dir;
    end
    if (sel) begin
      lineBuffer_511_value <= lineBuffer_510_value;
    end
    if (sel) begin
      lineBuffer_512_value <= lineBuffer_511_value;
    end
    if (sel) begin
      lineBuffer_513_value <= lineBuffer_512_value;
    end
    if (sel) begin
      lineBuffer_514_value <= lineBuffer_513_value;
    end
    if (sel) begin
      lineBuffer_515_value <= lineBuffer_514_value;
    end
    if (sel) begin
      lineBuffer_516_value <= lineBuffer_515_value;
    end
    if (sel) begin
      lineBuffer_517_value <= lineBuffer_516_value;
    end
    if (sel) begin
      lineBuffer_518_value <= lineBuffer_517_value;
    end
    if (sel) begin
      lineBuffer_519_value <= lineBuffer_518_value;
    end
    if (sel) begin
      lineBuffer_520_value <= lineBuffer_519_value;
    end
    if (sel) begin
      lineBuffer_521_value <= lineBuffer_520_value;
    end
    if (sel) begin
      lineBuffer_522_value <= lineBuffer_521_value;
    end
    if (sel) begin
      lineBuffer_523_value <= lineBuffer_522_value;
    end
    if (sel) begin
      lineBuffer_524_value <= lineBuffer_523_value;
    end
    if (sel) begin
      lineBuffer_525_value <= lineBuffer_524_value;
    end
    if (sel) begin
      lineBuffer_526_value <= lineBuffer_525_value;
    end
    if (sel) begin
      lineBuffer_527_value <= lineBuffer_526_value;
    end
    if (sel) begin
      lineBuffer_528_value <= lineBuffer_527_value;
    end
    if (sel) begin
      lineBuffer_529_value <= lineBuffer_528_value;
    end
    if (sel) begin
      lineBuffer_530_value <= lineBuffer_529_value;
    end
    if (sel) begin
      lineBuffer_531_value <= lineBuffer_530_value;
    end
    if (sel) begin
      lineBuffer_532_value <= lineBuffer_531_value;
    end
    if (sel) begin
      lineBuffer_533_value <= lineBuffer_532_value;
    end
    if (sel) begin
      lineBuffer_534_value <= lineBuffer_533_value;
    end
    if (sel) begin
      lineBuffer_535_value <= lineBuffer_534_value;
    end
    if (sel) begin
      lineBuffer_536_value <= lineBuffer_535_value;
    end
    if (sel) begin
      lineBuffer_537_value <= lineBuffer_536_value;
    end
    if (sel) begin
      lineBuffer_538_value <= lineBuffer_537_value;
    end
    if (sel) begin
      lineBuffer_539_value <= lineBuffer_538_value;
    end
    if (sel) begin
      lineBuffer_540_value <= lineBuffer_539_value;
    end
    if (sel) begin
      lineBuffer_541_value <= lineBuffer_540_value;
    end
    if (sel) begin
      lineBuffer_542_value <= lineBuffer_541_value;
    end
    if (sel) begin
      lineBuffer_543_value <= lineBuffer_542_value;
    end
    if (sel) begin
      lineBuffer_544_value <= lineBuffer_543_value;
    end
    if (sel) begin
      lineBuffer_545_value <= lineBuffer_544_value;
    end
    if (sel) begin
      lineBuffer_546_value <= lineBuffer_545_value;
    end
    if (sel) begin
      lineBuffer_547_value <= lineBuffer_546_value;
    end
    if (sel) begin
      lineBuffer_548_value <= lineBuffer_547_value;
    end
    if (sel) begin
      lineBuffer_549_value <= lineBuffer_548_value;
    end
    if (sel) begin
      lineBuffer_550_value <= lineBuffer_549_value;
    end
    if (sel) begin
      lineBuffer_551_value <= lineBuffer_550_value;
    end
    if (sel) begin
      lineBuffer_552_value <= lineBuffer_551_value;
    end
    if (sel) begin
      lineBuffer_553_value <= lineBuffer_552_value;
    end
    if (sel) begin
      lineBuffer_554_value <= lineBuffer_553_value;
    end
    if (sel) begin
      lineBuffer_555_value <= lineBuffer_554_value;
    end
    if (sel) begin
      lineBuffer_556_value <= lineBuffer_555_value;
    end
    if (sel) begin
      lineBuffer_557_value <= lineBuffer_556_value;
    end
    if (sel) begin
      lineBuffer_558_value <= lineBuffer_557_value;
    end
    if (sel) begin
      lineBuffer_559_value <= lineBuffer_558_value;
    end
    if (sel) begin
      lineBuffer_560_value <= lineBuffer_559_value;
    end
    if (sel) begin
      lineBuffer_561_value <= lineBuffer_560_value;
    end
    if (sel) begin
      lineBuffer_562_value <= lineBuffer_561_value;
    end
    if (sel) begin
      lineBuffer_563_value <= lineBuffer_562_value;
    end
    if (sel) begin
      lineBuffer_564_value <= lineBuffer_563_value;
    end
    if (sel) begin
      lineBuffer_565_value <= lineBuffer_564_value;
    end
    if (sel) begin
      lineBuffer_566_value <= lineBuffer_565_value;
    end
    if (sel) begin
      lineBuffer_567_value <= lineBuffer_566_value;
    end
    if (sel) begin
      lineBuffer_568_value <= lineBuffer_567_value;
    end
    if (sel) begin
      lineBuffer_569_value <= lineBuffer_568_value;
    end
    if (sel) begin
      lineBuffer_570_value <= lineBuffer_569_value;
    end
    if (sel) begin
      lineBuffer_571_value <= lineBuffer_570_value;
    end
    if (sel) begin
      lineBuffer_572_value <= lineBuffer_571_value;
    end
    if (sel) begin
      lineBuffer_573_value <= lineBuffer_572_value;
    end
    if (sel) begin
      lineBuffer_574_value <= lineBuffer_573_value;
    end
    if (sel) begin
      lineBuffer_575_value <= lineBuffer_574_value;
    end
    if (sel) begin
      lineBuffer_576_value <= lineBuffer_575_value;
    end
    if (sel) begin
      lineBuffer_577_value <= lineBuffer_576_value;
    end
    if (sel) begin
      lineBuffer_578_value <= lineBuffer_577_value;
    end
    if (sel) begin
      lineBuffer_579_value <= lineBuffer_578_value;
    end
    if (sel) begin
      lineBuffer_580_value <= lineBuffer_579_value;
    end
    if (sel) begin
      lineBuffer_581_value <= lineBuffer_580_value;
    end
    if (sel) begin
      lineBuffer_582_value <= lineBuffer_581_value;
    end
    if (sel) begin
      lineBuffer_583_value <= lineBuffer_582_value;
    end
    if (sel) begin
      lineBuffer_584_value <= lineBuffer_583_value;
    end
    if (sel) begin
      lineBuffer_585_value <= lineBuffer_584_value;
    end
    if (sel) begin
      lineBuffer_586_value <= lineBuffer_585_value;
    end
    if (sel) begin
      lineBuffer_587_value <= lineBuffer_586_value;
    end
    if (sel) begin
      lineBuffer_588_value <= lineBuffer_587_value;
    end
    if (sel) begin
      lineBuffer_589_value <= lineBuffer_588_value;
    end
    if (sel) begin
      lineBuffer_590_value <= lineBuffer_589_value;
    end
    if (sel) begin
      lineBuffer_591_value <= lineBuffer_590_value;
    end
    if (sel) begin
      lineBuffer_592_value <= lineBuffer_591_value;
    end
    if (sel) begin
      lineBuffer_593_value <= lineBuffer_592_value;
    end
    if (sel) begin
      lineBuffer_594_value <= lineBuffer_593_value;
    end
    if (sel) begin
      lineBuffer_595_value <= lineBuffer_594_value;
    end
    if (sel) begin
      lineBuffer_596_value <= lineBuffer_595_value;
    end
    if (sel) begin
      lineBuffer_597_value <= lineBuffer_596_value;
    end
    if (sel) begin
      lineBuffer_598_value <= lineBuffer_597_value;
    end
    if (sel) begin
      lineBuffer_599_value <= lineBuffer_598_value;
    end
    if (sel) begin
      lineBuffer_600_value <= lineBuffer_599_value;
    end
    if (sel) begin
      lineBuffer_601_value <= lineBuffer_600_value;
    end
    if (sel) begin
      lineBuffer_602_value <= lineBuffer_601_value;
    end
    if (sel) begin
      lineBuffer_603_value <= lineBuffer_602_value;
    end
    if (sel) begin
      lineBuffer_604_value <= lineBuffer_603_value;
    end
    if (sel) begin
      lineBuffer_605_value <= lineBuffer_604_value;
    end
    if (sel) begin
      lineBuffer_606_value <= lineBuffer_605_value;
    end
    if (sel) begin
      lineBuffer_607_value <= lineBuffer_606_value;
    end
    if (sel) begin
      lineBuffer_608_value <= lineBuffer_607_value;
    end
    if (sel) begin
      lineBuffer_609_value <= lineBuffer_608_value;
    end
    if (sel) begin
      lineBuffer_610_value <= lineBuffer_609_value;
    end
    if (sel) begin
      lineBuffer_611_value <= lineBuffer_610_value;
    end
    if (sel) begin
      lineBuffer_612_value <= lineBuffer_611_value;
    end
    if (sel) begin
      lineBuffer_613_value <= lineBuffer_612_value;
    end
    if (sel) begin
      lineBuffer_614_value <= lineBuffer_613_value;
    end
    if (sel) begin
      lineBuffer_615_value <= lineBuffer_614_value;
    end
    if (sel) begin
      lineBuffer_616_value <= lineBuffer_615_value;
    end
    if (sel) begin
      lineBuffer_617_value <= lineBuffer_616_value;
    end
    if (sel) begin
      lineBuffer_618_value <= lineBuffer_617_value;
    end
    if (sel) begin
      lineBuffer_619_value <= lineBuffer_618_value;
    end
    if (sel) begin
      lineBuffer_620_value <= lineBuffer_619_value;
    end
    if (sel) begin
      lineBuffer_621_value <= lineBuffer_620_value;
    end
    if (sel) begin
      lineBuffer_622_value <= lineBuffer_621_value;
    end
    if (sel) begin
      lineBuffer_623_value <= lineBuffer_622_value;
    end
    if (sel) begin
      lineBuffer_624_value <= lineBuffer_623_value;
    end
    if (sel) begin
      lineBuffer_625_value <= lineBuffer_624_value;
    end
    if (sel) begin
      lineBuffer_626_value <= lineBuffer_625_value;
    end
    if (sel) begin
      lineBuffer_627_value <= lineBuffer_626_value;
    end
    if (sel) begin
      lineBuffer_628_value <= lineBuffer_627_value;
    end
    if (sel) begin
      lineBuffer_629_value <= lineBuffer_628_value;
    end
    if (sel) begin
      lineBuffer_630_value <= lineBuffer_629_value;
    end
    if (sel) begin
      lineBuffer_631_value <= lineBuffer_630_value;
    end
    if (sel) begin
      lineBuffer_632_value <= lineBuffer_631_value;
    end
    if (sel) begin
      lineBuffer_633_value <= lineBuffer_632_value;
    end
    if (sel) begin
      lineBuffer_634_value <= lineBuffer_633_value;
    end
    if (sel) begin
      lineBuffer_635_value <= lineBuffer_634_value;
    end
    if (sel) begin
      lineBuffer_636_value <= lineBuffer_635_value;
    end
    if (sel) begin
      lineBuffer_637_value <= lineBuffer_636_value;
    end
    if (sel) begin
      lineBuffer_638_value <= lineBuffer_637_value;
    end
    if (sel) begin
      lineBuffer_639_value <= lineBuffer_638_value;
    end
    if (sel) begin
      lineBuffer_640_value <= lineBuffer_639_value;
    end
    if (sel) begin
      lineBuffer_641_value <= lineBuffer_640_value;
    end
    if (sel) begin
      lineBuffer_642_value <= lineBuffer_641_value;
    end
    if (sel) begin
      lineBuffer_643_value <= lineBuffer_642_value;
    end
    if (sel) begin
      lineBuffer_644_value <= lineBuffer_643_value;
    end
    if (sel) begin
      lineBuffer_645_value <= lineBuffer_644_value;
    end
    if (sel) begin
      lineBuffer_646_value <= lineBuffer_645_value;
    end
    if (sel) begin
      lineBuffer_647_value <= lineBuffer_646_value;
    end
    if (sel) begin
      lineBuffer_648_value <= lineBuffer_647_value;
    end
    if (sel) begin
      lineBuffer_649_value <= lineBuffer_648_value;
    end
    if (sel) begin
      lineBuffer_650_value <= lineBuffer_649_value;
    end
    if (sel) begin
      lineBuffer_651_value <= lineBuffer_650_value;
    end
    if (sel) begin
      lineBuffer_652_value <= lineBuffer_651_value;
    end
    if (sel) begin
      lineBuffer_653_value <= lineBuffer_652_value;
    end
    if (sel) begin
      lineBuffer_654_value <= lineBuffer_653_value;
    end
    if (sel) begin
      lineBuffer_655_value <= lineBuffer_654_value;
    end
    if (sel) begin
      lineBuffer_656_value <= lineBuffer_655_value;
    end
    if (sel) begin
      lineBuffer_657_value <= lineBuffer_656_value;
    end
    if (sel) begin
      lineBuffer_658_value <= lineBuffer_657_value;
    end
    if (sel) begin
      lineBuffer_659_value <= lineBuffer_658_value;
    end
    if (sel) begin
      lineBuffer_660_value <= lineBuffer_659_value;
    end
    if (sel) begin
      lineBuffer_661_value <= lineBuffer_660_value;
    end
    if (sel) begin
      lineBuffer_662_value <= lineBuffer_661_value;
    end
    if (sel) begin
      lineBuffer_663_value <= lineBuffer_662_value;
    end
    if (sel) begin
      lineBuffer_664_value <= lineBuffer_663_value;
    end
    if (sel) begin
      lineBuffer_665_value <= lineBuffer_664_value;
    end
    if (sel) begin
      lineBuffer_666_value <= lineBuffer_665_value;
    end
    if (sel) begin
      lineBuffer_667_value <= lineBuffer_666_value;
    end
    if (sel) begin
      lineBuffer_668_value <= lineBuffer_667_value;
    end
    if (sel) begin
      lineBuffer_669_value <= lineBuffer_668_value;
    end
    if (sel) begin
      lineBuffer_670_value <= lineBuffer_669_value;
    end
    if (sel) begin
      lineBuffer_671_value <= lineBuffer_670_value;
    end
    if (sel) begin
      lineBuffer_672_value <= lineBuffer_671_value;
    end
    if (sel) begin
      lineBuffer_673_value <= lineBuffer_672_value;
    end
    if (sel) begin
      lineBuffer_674_value <= lineBuffer_673_value;
    end
    if (sel) begin
      lineBuffer_675_value <= lineBuffer_674_value;
    end
    if (sel) begin
      lineBuffer_676_value <= lineBuffer_675_value;
    end
    if (sel) begin
      lineBuffer_677_value <= lineBuffer_676_value;
    end
    if (sel) begin
      lineBuffer_678_value <= lineBuffer_677_value;
    end
    if (sel) begin
      lineBuffer_679_value <= lineBuffer_678_value;
    end
    if (sel) begin
      lineBuffer_680_value <= lineBuffer_679_value;
    end
    if (sel) begin
      lineBuffer_681_value <= lineBuffer_680_value;
    end
    if (sel) begin
      lineBuffer_682_value <= lineBuffer_681_value;
    end
    if (sel) begin
      lineBuffer_683_value <= lineBuffer_682_value;
    end
    if (sel) begin
      lineBuffer_684_value <= lineBuffer_683_value;
    end
    if (sel) begin
      lineBuffer_685_value <= lineBuffer_684_value;
    end
    if (sel) begin
      lineBuffer_686_value <= lineBuffer_685_value;
    end
    if (sel) begin
      lineBuffer_687_value <= lineBuffer_686_value;
    end
    if (sel) begin
      lineBuffer_688_value <= lineBuffer_687_value;
    end
    if (sel) begin
      lineBuffer_689_value <= lineBuffer_688_value;
    end
    if (sel) begin
      lineBuffer_690_value <= lineBuffer_689_value;
    end
    if (sel) begin
      lineBuffer_691_value <= lineBuffer_690_value;
    end
    if (sel) begin
      lineBuffer_692_value <= lineBuffer_691_value;
    end
    if (sel) begin
      lineBuffer_693_value <= lineBuffer_692_value;
    end
    if (sel) begin
      lineBuffer_694_value <= lineBuffer_693_value;
    end
    if (sel) begin
      lineBuffer_695_value <= lineBuffer_694_value;
    end
    if (sel) begin
      lineBuffer_696_value <= lineBuffer_695_value;
    end
    if (sel) begin
      lineBuffer_697_value <= lineBuffer_696_value;
    end
    if (sel) begin
      lineBuffer_698_value <= lineBuffer_697_value;
    end
    if (sel) begin
      lineBuffer_699_value <= lineBuffer_698_value;
    end
    if (sel) begin
      lineBuffer_700_value <= lineBuffer_699_value;
    end
    if (sel) begin
      lineBuffer_701_value <= lineBuffer_700_value;
    end
    if (sel) begin
      lineBuffer_702_value <= lineBuffer_701_value;
    end
    if (sel) begin
      lineBuffer_703_value <= lineBuffer_702_value;
    end
    if (sel) begin
      lineBuffer_704_value <= lineBuffer_703_value;
    end
    if (sel) begin
      lineBuffer_705_value <= lineBuffer_704_value;
    end
    if (sel) begin
      lineBuffer_706_value <= lineBuffer_705_value;
    end
    if (sel) begin
      lineBuffer_707_value <= lineBuffer_706_value;
    end
    if (sel) begin
      lineBuffer_708_value <= lineBuffer_707_value;
    end
    if (sel) begin
      lineBuffer_709_value <= lineBuffer_708_value;
    end
    if (sel) begin
      lineBuffer_710_value <= lineBuffer_709_value;
    end
    if (sel) begin
      lineBuffer_711_value <= lineBuffer_710_value;
    end
    if (sel) begin
      lineBuffer_712_value <= lineBuffer_711_value;
    end
    if (sel) begin
      lineBuffer_713_value <= lineBuffer_712_value;
    end
    if (sel) begin
      lineBuffer_714_value <= lineBuffer_713_value;
    end
    if (sel) begin
      lineBuffer_715_value <= lineBuffer_714_value;
    end
    if (sel) begin
      lineBuffer_716_value <= lineBuffer_715_value;
    end
    if (sel) begin
      lineBuffer_717_value <= lineBuffer_716_value;
    end
    if (sel) begin
      lineBuffer_718_value <= lineBuffer_717_value;
    end
    if (sel) begin
      lineBuffer_719_value <= lineBuffer_718_value;
    end
    if (sel) begin
      lineBuffer_720_value <= lineBuffer_719_value;
    end
    if (sel) begin
      lineBuffer_721_value <= lineBuffer_720_value;
    end
    if (sel) begin
      lineBuffer_722_value <= lineBuffer_721_value;
    end
    if (sel) begin
      lineBuffer_723_value <= lineBuffer_722_value;
    end
    if (sel) begin
      lineBuffer_724_value <= lineBuffer_723_value;
    end
    if (sel) begin
      lineBuffer_725_value <= lineBuffer_724_value;
    end
    if (sel) begin
      lineBuffer_726_value <= lineBuffer_725_value;
    end
    if (sel) begin
      lineBuffer_727_value <= lineBuffer_726_value;
    end
    if (sel) begin
      lineBuffer_728_value <= lineBuffer_727_value;
    end
    if (sel) begin
      lineBuffer_729_value <= lineBuffer_728_value;
    end
    if (sel) begin
      lineBuffer_730_value <= lineBuffer_729_value;
    end
    if (sel) begin
      lineBuffer_731_value <= lineBuffer_730_value;
    end
    if (sel) begin
      lineBuffer_732_value <= lineBuffer_731_value;
    end
    if (sel) begin
      lineBuffer_733_value <= lineBuffer_732_value;
    end
    if (sel) begin
      lineBuffer_734_value <= lineBuffer_733_value;
    end
    if (sel) begin
      lineBuffer_735_value <= lineBuffer_734_value;
    end
    if (sel) begin
      lineBuffer_736_value <= lineBuffer_735_value;
    end
    if (sel) begin
      lineBuffer_737_value <= lineBuffer_736_value;
    end
    if (sel) begin
      lineBuffer_738_value <= lineBuffer_737_value;
    end
    if (sel) begin
      lineBuffer_739_value <= lineBuffer_738_value;
    end
    if (sel) begin
      lineBuffer_740_value <= lineBuffer_739_value;
    end
    if (sel) begin
      lineBuffer_741_value <= lineBuffer_740_value;
    end
    if (sel) begin
      lineBuffer_742_value <= lineBuffer_741_value;
    end
    if (sel) begin
      lineBuffer_743_value <= lineBuffer_742_value;
    end
    if (sel) begin
      lineBuffer_744_value <= lineBuffer_743_value;
    end
    if (sel) begin
      lineBuffer_745_value <= lineBuffer_744_value;
    end
    if (sel) begin
      lineBuffer_746_value <= lineBuffer_745_value;
    end
    if (sel) begin
      lineBuffer_747_value <= lineBuffer_746_value;
    end
    if (sel) begin
      lineBuffer_748_value <= lineBuffer_747_value;
    end
    if (sel) begin
      lineBuffer_749_value <= lineBuffer_748_value;
    end
    if (sel) begin
      lineBuffer_750_value <= lineBuffer_749_value;
    end
    if (sel) begin
      lineBuffer_751_value <= lineBuffer_750_value;
    end
    if (sel) begin
      lineBuffer_752_value <= lineBuffer_751_value;
    end
    if (sel) begin
      lineBuffer_753_value <= lineBuffer_752_value;
    end
    if (sel) begin
      lineBuffer_754_value <= lineBuffer_753_value;
    end
    if (sel) begin
      lineBuffer_755_value <= lineBuffer_754_value;
    end
    if (sel) begin
      lineBuffer_756_value <= lineBuffer_755_value;
    end
    if (sel) begin
      lineBuffer_757_value <= lineBuffer_756_value;
    end
    if (sel) begin
      lineBuffer_758_value <= lineBuffer_757_value;
    end
    if (sel) begin
      lineBuffer_759_value <= lineBuffer_758_value;
    end
    if (sel) begin
      lineBuffer_760_value <= lineBuffer_759_value;
    end
    if (sel) begin
      lineBuffer_761_value <= lineBuffer_760_value;
    end
    if (sel) begin
      lineBuffer_762_value <= lineBuffer_761_value;
    end
    if (sel) begin
      lineBuffer_763_value <= lineBuffer_762_value;
    end
    if (sel) begin
      lineBuffer_764_value <= lineBuffer_763_value;
    end
    if (sel) begin
      lineBuffer_765_value <= lineBuffer_764_value;
    end
    if (sel) begin
      lineBuffer_766_value <= lineBuffer_765_value;
    end
    if (sel) begin
      lineBuffer_767_value <= lineBuffer_766_value;
    end
    if (sel) begin
      windowBuffer_0_value <= windowBuffer_1_value;
    end
    if (sel) begin
      windowBuffer_1_value <= windowBuffer_2_value;
    end
    if (sel) begin
      windowBuffer_2_value <= lineBuffer_255_value;
    end
    if (sel) begin
      windowBuffer_3_value <= windowBuffer_4_value;
    end
    if (sel) begin
      windowBuffer_4_grad_dir <= windowBuffer_5_grad_dir;
    end
    if (sel) begin
      windowBuffer_4_value <= windowBuffer_5_value;
    end
    if (sel) begin
      windowBuffer_5_grad_dir <= lineBuffer_511_grad_dir;
    end
    if (sel) begin
      windowBuffer_5_value <= lineBuffer_511_value;
    end
    if (sel) begin
      windowBuffer_6_value <= windowBuffer_7_value;
    end
    if (sel) begin
      windowBuffer_7_value <= windowBuffer_8_value;
    end
    if (sel) begin
      windowBuffer_8_value <= lineBuffer_767_value;
    end
  end
endmodule
module SobelAndNonMaxSupressionFilter(
  input        clock,
  input        reset,
  output       io_enq_ready,
  input        io_enq_valid,
  input  [7:0] io_enq_bits,
  input        io_enq_user,
  input        io_enq_last,
  input        io_deq_ready,
  output       io_deq_valid,
  output [7:0] io_deq_bits,
  output       io_deq_user,
  output       io_deq_last
);
  wire  sobel_clock; // @[ChiselImProc.scala 411:24]
  wire  sobel_reset; // @[ChiselImProc.scala 411:24]
  wire  sobel_io_enq_ready; // @[ChiselImProc.scala 411:24]
  wire  sobel_io_enq_valid; // @[ChiselImProc.scala 411:24]
  wire [7:0] sobel_io_enq_bits; // @[ChiselImProc.scala 411:24]
  wire  sobel_io_enq_user; // @[ChiselImProc.scala 411:24]
  wire  sobel_io_enq_last; // @[ChiselImProc.scala 411:24]
  wire  sobel_io_deq_ready; // @[ChiselImProc.scala 411:24]
  wire  sobel_io_deq_valid; // @[ChiselImProc.scala 411:24]
  wire [1:0] sobel_io_deq_bits_grad_dir; // @[ChiselImProc.scala 411:24]
  wire [7:0] sobel_io_deq_bits_value; // @[ChiselImProc.scala 411:24]
  wire  sobel_io_deq_user; // @[ChiselImProc.scala 411:24]
  wire  sobel_io_deq_last; // @[ChiselImProc.scala 411:24]
  wire  nonmaxSupression_clock; // @[ChiselImProc.scala 412:35]
  wire  nonmaxSupression_reset; // @[ChiselImProc.scala 412:35]
  wire  nonmaxSupression_io_enq_ready; // @[ChiselImProc.scala 412:35]
  wire  nonmaxSupression_io_enq_valid; // @[ChiselImProc.scala 412:35]
  wire [1:0] nonmaxSupression_io_enq_bits_grad_dir; // @[ChiselImProc.scala 412:35]
  wire [7:0] nonmaxSupression_io_enq_bits_value; // @[ChiselImProc.scala 412:35]
  wire  nonmaxSupression_io_enq_user; // @[ChiselImProc.scala 412:35]
  wire  nonmaxSupression_io_enq_last; // @[ChiselImProc.scala 412:35]
  wire  nonmaxSupression_io_deq_ready; // @[ChiselImProc.scala 412:35]
  wire  nonmaxSupression_io_deq_valid; // @[ChiselImProc.scala 412:35]
  wire [7:0] nonmaxSupression_io_deq_bits; // @[ChiselImProc.scala 412:35]
  wire  nonmaxSupression_io_deq_user; // @[ChiselImProc.scala 412:35]
  wire  nonmaxSupression_io_deq_last; // @[ChiselImProc.scala 412:35]
  SobelFilter sobel ( // @[ChiselImProc.scala 411:24]
    .clock(sobel_clock),
    .reset(sobel_reset),
    .io_enq_ready(sobel_io_enq_ready),
    .io_enq_valid(sobel_io_enq_valid),
    .io_enq_bits(sobel_io_enq_bits),
    .io_enq_user(sobel_io_enq_user),
    .io_enq_last(sobel_io_enq_last),
    .io_deq_ready(sobel_io_deq_ready),
    .io_deq_valid(sobel_io_deq_valid),
    .io_deq_bits_grad_dir(sobel_io_deq_bits_grad_dir),
    .io_deq_bits_value(sobel_io_deq_bits_value),
    .io_deq_user(sobel_io_deq_user),
    .io_deq_last(sobel_io_deq_last)
  );
  NonMaxSupression nonmaxSupression ( // @[ChiselImProc.scala 412:35]
    .clock(nonmaxSupression_clock),
    .reset(nonmaxSupression_reset),
    .io_enq_ready(nonmaxSupression_io_enq_ready),
    .io_enq_valid(nonmaxSupression_io_enq_valid),
    .io_enq_bits_grad_dir(nonmaxSupression_io_enq_bits_grad_dir),
    .io_enq_bits_value(nonmaxSupression_io_enq_bits_value),
    .io_enq_user(nonmaxSupression_io_enq_user),
    .io_enq_last(nonmaxSupression_io_enq_last),
    .io_deq_ready(nonmaxSupression_io_deq_ready),
    .io_deq_valid(nonmaxSupression_io_deq_valid),
    .io_deq_bits(nonmaxSupression_io_deq_bits),
    .io_deq_user(nonmaxSupression_io_deq_user),
    .io_deq_last(nonmaxSupression_io_deq_last)
  );
  assign io_enq_ready = sobel_io_enq_ready; // @[ChiselImProc.scala 116:22 ChiselImProc.scala 414:12]
  assign io_deq_valid = nonmaxSupression_io_deq_valid; // @[ChiselImProc.scala 117:22 ChiselImProc.scala 416:29]
  assign io_deq_bits = nonmaxSupression_io_deq_bits; // @[ChiselImProc.scala 416:29]
  assign io_deq_user = nonmaxSupression_io_deq_user; // @[ChiselImProc.scala 144:17 ChiselImProc.scala 114:21 ChiselImProc.scala 416:29]
  assign io_deq_last = nonmaxSupression_io_deq_last; // @[ChiselImProc.scala 143:17 ChiselImProc.scala 113:21 ChiselImProc.scala 416:29]
  assign sobel_clock = clock;
  assign sobel_reset = reset;
  assign sobel_io_enq_valid = io_enq_valid; // @[ChiselImProc.scala 414:12]
  assign sobel_io_enq_bits = io_enq_bits; // @[ChiselImProc.scala 414:12]
  assign sobel_io_enq_user = io_enq_user; // @[ChiselImProc.scala 414:12]
  assign sobel_io_enq_last = io_enq_last; // @[ChiselImProc.scala 414:12]
  assign sobel_io_deq_ready = nonmaxSupression_io_enq_ready; // @[ChiselImProc.scala 415:18]
  assign nonmaxSupression_clock = clock;
  assign nonmaxSupression_reset = reset;
  assign nonmaxSupression_io_enq_valid = sobel_io_deq_valid; // @[ChiselImProc.scala 415:18]
  assign nonmaxSupression_io_enq_bits_grad_dir = sobel_io_deq_bits_grad_dir; // @[ChiselImProc.scala 415:18]
  assign nonmaxSupression_io_enq_bits_value = sobel_io_deq_bits_value; // @[ChiselImProc.scala 415:18]
  assign nonmaxSupression_io_enq_user = sobel_io_deq_user; // @[ChiselImProc.scala 415:18]
  assign nonmaxSupression_io_enq_last = sobel_io_deq_last; // @[ChiselImProc.scala 415:18]
  assign nonmaxSupression_io_deq_ready = io_deq_ready; // @[ChiselImProc.scala 416:29]
endmodule
module ZeroPadding(
  input        clock,
  input        reset,
  output       io_enq_ready,
  input        io_enq_valid,
  input  [7:0] io_enq_bits,
  input        io_enq_user,
  input        io_enq_last,
  input        io_deq_ready,
  output       io_deq_valid,
  output [7:0] io_deq_bits,
  output       io_deq_user,
  output       io_deq_last
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
`endif // RANDOMIZE_REG_INIT
  reg [1:0] stateReg; // @[ChiselImProc.scala 62:28]
  reg [7:0] dataReg; // @[ChiselImProc.scala 64:23]
  reg [7:0] shadowReg; // @[ChiselImProc.scala 66:25]
  reg  userReg; // @[ChiselImProc.scala 67:23]
  reg  shadowUserReg; // @[ChiselImProc.scala 68:29]
  reg  lastReg; // @[ChiselImProc.scala 69:23]
  reg  shadowLastReg; // @[ChiselImProc.scala 70:29]
  wire  _T = 2'h0 == stateReg; // @[Conditional.scala 37:30]
  wire  _T_1 = 2'h1 == stateReg; // @[Conditional.scala 37:30]
  wire  _T_2 = ~io_enq_valid; // @[ChiselImProc.scala 84:39]
  wire  _T_3 = io_deq_ready & _T_2; // @[ChiselImProc.scala 84:36]
  wire  _T_4 = io_deq_ready & io_enq_valid; // @[ChiselImProc.scala 87:42]
  wire  _T_5 = ~io_deq_ready; // @[ChiselImProc.scala 92:29]
  wire  _T_6 = _T_5 & io_enq_valid; // @[ChiselImProc.scala 92:43]
  wire  _T_7 = 2'h2 == stateReg; // @[Conditional.scala 37:30]
  wire  _T_8 = 2'h3 == stateReg; // @[Conditional.scala 37:30]
  wire  _T_9 = stateReg == 2'h0; // @[ChiselImProc.scala 116:35]
  wire  _T_10 = stateReg == 2'h1; // @[ChiselImProc.scala 116:57]
  wire  _T_11 = _T_9 | _T_10; // @[ChiselImProc.scala 116:45]
  wire  _T_12 = stateReg == 2'h3; // @[ChiselImProc.scala 116:77]
  wire  _T_15 = stateReg == 2'h2; // @[ChiselImProc.scala 117:55]
  wire  _T_16 = _T_10 | _T_15; // @[ChiselImProc.scala 117:43]
  reg [8:0] xcounter; // @[ChiselImProc.scala 423:23]
  reg [8:0] ycounter; // @[ChiselImProc.scala 424:23]
  wire  _T_20 = lastReg & _T_16; // @[ChiselImProc.scala 429:25]
  wire  _T_21 = _T_20 & io_deq_ready; // @[ChiselImProc.scala 429:67]
  wire [8:0] _T_23 = ycounter + 9'h1; // @[ChiselImProc.scala 431:30]
  wire  _T_27 = _T_16 & io_deq_ready; // @[ChiselImProc.scala 432:56]
  wire [8:0] _T_29 = xcounter + 9'h1; // @[ChiselImProc.scala 433:30]
  wire  _T_30 = 9'h5 < xcounter; // @[ChiselImProc.scala 436:24]
  wire [8:0] _T_32 = 9'h100 - 9'h5; // @[ChiselImProc.scala 436:56]
  wire  _T_33 = xcounter < _T_32; // @[ChiselImProc.scala 436:47]
  wire  _T_34 = _T_30 & _T_33; // @[ChiselImProc.scala 436:35]
  wire  _T_35 = 9'h5 < ycounter; // @[ChiselImProc.scala 437:26]
  wire  _T_36 = _T_34 & _T_35; // @[ChiselImProc.scala 436:70]
  wire  _T_39 = ycounter < _T_32; // @[ChiselImProc.scala 437:49]
  wire  _T_40 = _T_36 & _T_39; // @[ChiselImProc.scala 437:37]
  assign io_enq_ready = _T_11 | _T_12; // @[ChiselImProc.scala 116:22]
  assign io_deq_valid = _T_10 | _T_15; // @[ChiselImProc.scala 117:22]
  assign io_deq_bits = _T_40 ? dataReg : 8'h0; // @[ChiselImProc.scala 438:21 ChiselImProc.scala 440:21]
  assign io_deq_user = userReg; // @[ChiselImProc.scala 144:17 ChiselImProc.scala 114:21]
  assign io_deq_last = lastReg; // @[ChiselImProc.scala 143:17 ChiselImProc.scala 113:21]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  stateReg = _RAND_0[1:0];
  _RAND_1 = {1{`RANDOM}};
  dataReg = _RAND_1[7:0];
  _RAND_2 = {1{`RANDOM}};
  shadowReg = _RAND_2[7:0];
  _RAND_3 = {1{`RANDOM}};
  userReg = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  shadowUserReg = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  lastReg = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  shadowLastReg = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  xcounter = _RAND_7[8:0];
  _RAND_8 = {1{`RANDOM}};
  ycounter = _RAND_8[8:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      stateReg <= 2'h0;
    end else if (_T) begin
      if (io_enq_valid) begin
        stateReg <= 2'h1;
      end
    end else if (_T_1) begin
      if (_T_3) begin
        stateReg <= 2'h0;
      end else if (_T_4) begin
        stateReg <= 2'h1;
      end else if (_T_6) begin
        stateReg <= 2'h2;
      end
    end else if (_T_7) begin
      if (io_deq_ready) begin
        stateReg <= 2'h1;
      end
    end else if (_T_8) begin
      stateReg <= 2'h0;
    end
    if (_T) begin
      if (io_enq_valid) begin
        dataReg <= io_enq_bits;
      end
    end else if (_T_1) begin
      if (!(_T_3)) begin
        if (_T_4) begin
          dataReg <= io_enq_bits;
        end
      end
    end else if (_T_7) begin
      if (io_deq_ready) begin
        dataReg <= shadowReg;
      end
    end
    if (!(_T)) begin
      if (_T_1) begin
        if (!(_T_3)) begin
          if (!(_T_4)) begin
            if (_T_6) begin
              shadowReg <= io_enq_bits;
            end
          end
        end
      end
    end
    if (_T) begin
      userReg <= io_enq_user;
    end else if (_T_1) begin
      if (_T_3) begin
        userReg <= io_enq_user;
      end else if (_T_4) begin
        userReg <= io_enq_user;
      end
    end else if (_T_7) begin
      if (io_deq_ready) begin
        userReg <= shadowUserReg;
      end
    end
    if (!(_T)) begin
      if (_T_1) begin
        if (!(_T_3)) begin
          if (!(_T_4)) begin
            if (_T_6) begin
              shadowUserReg <= io_enq_user;
            end
          end
        end
      end
    end
    if (_T) begin
      if (io_enq_valid) begin
        lastReg <= io_enq_last;
      end
    end else if (_T_1) begin
      if (!(_T_3)) begin
        if (_T_4) begin
          lastReg <= io_enq_last;
        end
      end
    end else if (_T_7) begin
      if (io_deq_ready) begin
        lastReg <= shadowLastReg;
      end
    end
    if (!(_T)) begin
      if (_T_1) begin
        if (!(_T_3)) begin
          if (!(_T_4)) begin
            if (_T_6) begin
              shadowLastReg <= io_enq_last;
            end
          end
        end
      end
    end
    if (userReg) begin
      xcounter <= 9'h0;
    end else if (_T_21) begin
      xcounter <= 9'h0;
    end else if (_T_27) begin
      xcounter <= _T_29;
    end
    if (userReg) begin
      ycounter <= 9'h0;
    end else if (_T_21) begin
      ycounter <= _T_23;
    end
  end
endmodule
module HystThreshold(
  input        clock,
  input        reset,
  output       io_enq_ready,
  input        io_enq_valid,
  input  [7:0] io_enq_bits,
  input        io_enq_user,
  input        io_enq_last,
  input        io_deq_ready,
  output       io_deq_valid,
  output [7:0] io_deq_bits,
  output       io_deq_user,
  output       io_deq_last
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
`endif // RANDOMIZE_REG_INIT
  reg [1:0] stateReg; // @[ChiselImProc.scala 62:28]
  reg [7:0] dataReg; // @[ChiselImProc.scala 64:23]
  reg [7:0] shadowReg; // @[ChiselImProc.scala 66:25]
  reg  userReg; // @[ChiselImProc.scala 67:23]
  reg  shadowUserReg; // @[ChiselImProc.scala 68:29]
  reg  lastReg; // @[ChiselImProc.scala 69:23]
  reg  shadowLastReg; // @[ChiselImProc.scala 70:29]
  wire  _T = 2'h0 == stateReg; // @[Conditional.scala 37:30]
  wire  _T_1 = 2'h1 == stateReg; // @[Conditional.scala 37:30]
  wire  _T_2 = ~io_enq_valid; // @[ChiselImProc.scala 84:39]
  wire  _T_3 = io_deq_ready & _T_2; // @[ChiselImProc.scala 84:36]
  wire  _T_4 = io_deq_ready & io_enq_valid; // @[ChiselImProc.scala 87:42]
  wire  _T_5 = ~io_deq_ready; // @[ChiselImProc.scala 92:29]
  wire  _T_6 = _T_5 & io_enq_valid; // @[ChiselImProc.scala 92:43]
  wire  _T_7 = 2'h2 == stateReg; // @[Conditional.scala 37:30]
  wire  _T_8 = 2'h3 == stateReg; // @[Conditional.scala 37:30]
  wire  _T_9 = stateReg == 2'h0; // @[ChiselImProc.scala 116:35]
  wire  _T_10 = stateReg == 2'h1; // @[ChiselImProc.scala 116:57]
  wire  _T_11 = _T_9 | _T_10; // @[ChiselImProc.scala 116:45]
  wire  _T_12 = stateReg == 2'h3; // @[ChiselImProc.scala 116:77]
  wire  _T_15 = stateReg == 2'h2; // @[ChiselImProc.scala 117:55]
  wire  _T_17 = dataReg < 8'h14; // @[ChiselImProc.scala 448:19]
  wire  _T_18 = dataReg > 8'h50; // @[ChiselImProc.scala 450:25]
  wire [7:0] _GEN_44 = _T_18 ? 8'hff : 8'h1; // @[ChiselImProc.scala 450:33]
  assign io_enq_ready = _T_11 | _T_12; // @[ChiselImProc.scala 116:22]
  assign io_deq_valid = _T_10 | _T_15; // @[ChiselImProc.scala 117:22]
  assign io_deq_bits = _T_17 ? 8'h0 : _GEN_44; // @[ChiselImProc.scala 449:21 ChiselImProc.scala 451:21 ChiselImProc.scala 453:21]
  assign io_deq_user = userReg; // @[ChiselImProc.scala 144:17 ChiselImProc.scala 114:21]
  assign io_deq_last = lastReg; // @[ChiselImProc.scala 143:17 ChiselImProc.scala 113:21]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  stateReg = _RAND_0[1:0];
  _RAND_1 = {1{`RANDOM}};
  dataReg = _RAND_1[7:0];
  _RAND_2 = {1{`RANDOM}};
  shadowReg = _RAND_2[7:0];
  _RAND_3 = {1{`RANDOM}};
  userReg = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  shadowUserReg = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  lastReg = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  shadowLastReg = _RAND_6[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      stateReg <= 2'h0;
    end else if (_T) begin
      if (io_enq_valid) begin
        stateReg <= 2'h1;
      end
    end else if (_T_1) begin
      if (_T_3) begin
        stateReg <= 2'h0;
      end else if (_T_4) begin
        stateReg <= 2'h1;
      end else if (_T_6) begin
        stateReg <= 2'h2;
      end
    end else if (_T_7) begin
      if (io_deq_ready) begin
        stateReg <= 2'h1;
      end
    end else if (_T_8) begin
      stateReg <= 2'h0;
    end
    if (_T) begin
      if (io_enq_valid) begin
        dataReg <= io_enq_bits;
      end
    end else if (_T_1) begin
      if (!(_T_3)) begin
        if (_T_4) begin
          dataReg <= io_enq_bits;
        end
      end
    end else if (_T_7) begin
      if (io_deq_ready) begin
        dataReg <= shadowReg;
      end
    end
    if (!(_T)) begin
      if (_T_1) begin
        if (!(_T_3)) begin
          if (!(_T_4)) begin
            if (_T_6) begin
              shadowReg <= io_enq_bits;
            end
          end
        end
      end
    end
    if (_T) begin
      userReg <= io_enq_user;
    end else if (_T_1) begin
      if (_T_3) begin
        userReg <= io_enq_user;
      end else if (_T_4) begin
        userReg <= io_enq_user;
      end
    end else if (_T_7) begin
      if (io_deq_ready) begin
        userReg <= shadowUserReg;
      end
    end
    if (!(_T)) begin
      if (_T_1) begin
        if (!(_T_3)) begin
          if (!(_T_4)) begin
            if (_T_6) begin
              shadowUserReg <= io_enq_user;
            end
          end
        end
      end
    end
    if (_T) begin
      if (io_enq_valid) begin
        lastReg <= io_enq_last;
      end
    end else if (_T_1) begin
      if (!(_T_3)) begin
        if (_T_4) begin
          lastReg <= io_enq_last;
        end
      end
    end else if (_T_7) begin
      if (io_deq_ready) begin
        lastReg <= shadowLastReg;
      end
    end
    if (!(_T)) begin
      if (_T_1) begin
        if (!(_T_3)) begin
          if (!(_T_4)) begin
            if (_T_6) begin
              shadowLastReg <= io_enq_last;
            end
          end
        end
      end
    end
  end
endmodule
module HystThresholdComp(
  input        clock,
  input        reset,
  output       io_enq_ready,
  input        io_enq_valid,
  input  [7:0] io_enq_bits,
  input        io_enq_user,
  input        io_enq_last,
  input        io_deq_ready,
  output       io_deq_valid,
  output [7:0] io_deq_bits,
  output       io_deq_user,
  output       io_deq_last
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
  reg [31:0] _RAND_64;
  reg [31:0] _RAND_65;
  reg [31:0] _RAND_66;
  reg [31:0] _RAND_67;
  reg [31:0] _RAND_68;
  reg [31:0] _RAND_69;
  reg [31:0] _RAND_70;
  reg [31:0] _RAND_71;
  reg [31:0] _RAND_72;
  reg [31:0] _RAND_73;
  reg [31:0] _RAND_74;
  reg [31:0] _RAND_75;
  reg [31:0] _RAND_76;
  reg [31:0] _RAND_77;
  reg [31:0] _RAND_78;
  reg [31:0] _RAND_79;
  reg [31:0] _RAND_80;
  reg [31:0] _RAND_81;
  reg [31:0] _RAND_82;
  reg [31:0] _RAND_83;
  reg [31:0] _RAND_84;
  reg [31:0] _RAND_85;
  reg [31:0] _RAND_86;
  reg [31:0] _RAND_87;
  reg [31:0] _RAND_88;
  reg [31:0] _RAND_89;
  reg [31:0] _RAND_90;
  reg [31:0] _RAND_91;
  reg [31:0] _RAND_92;
  reg [31:0] _RAND_93;
  reg [31:0] _RAND_94;
  reg [31:0] _RAND_95;
  reg [31:0] _RAND_96;
  reg [31:0] _RAND_97;
  reg [31:0] _RAND_98;
  reg [31:0] _RAND_99;
  reg [31:0] _RAND_100;
  reg [31:0] _RAND_101;
  reg [31:0] _RAND_102;
  reg [31:0] _RAND_103;
  reg [31:0] _RAND_104;
  reg [31:0] _RAND_105;
  reg [31:0] _RAND_106;
  reg [31:0] _RAND_107;
  reg [31:0] _RAND_108;
  reg [31:0] _RAND_109;
  reg [31:0] _RAND_110;
  reg [31:0] _RAND_111;
  reg [31:0] _RAND_112;
  reg [31:0] _RAND_113;
  reg [31:0] _RAND_114;
  reg [31:0] _RAND_115;
  reg [31:0] _RAND_116;
  reg [31:0] _RAND_117;
  reg [31:0] _RAND_118;
  reg [31:0] _RAND_119;
  reg [31:0] _RAND_120;
  reg [31:0] _RAND_121;
  reg [31:0] _RAND_122;
  reg [31:0] _RAND_123;
  reg [31:0] _RAND_124;
  reg [31:0] _RAND_125;
  reg [31:0] _RAND_126;
  reg [31:0] _RAND_127;
  reg [31:0] _RAND_128;
  reg [31:0] _RAND_129;
  reg [31:0] _RAND_130;
  reg [31:0] _RAND_131;
  reg [31:0] _RAND_132;
  reg [31:0] _RAND_133;
  reg [31:0] _RAND_134;
  reg [31:0] _RAND_135;
  reg [31:0] _RAND_136;
  reg [31:0] _RAND_137;
  reg [31:0] _RAND_138;
  reg [31:0] _RAND_139;
  reg [31:0] _RAND_140;
  reg [31:0] _RAND_141;
  reg [31:0] _RAND_142;
  reg [31:0] _RAND_143;
  reg [31:0] _RAND_144;
  reg [31:0] _RAND_145;
  reg [31:0] _RAND_146;
  reg [31:0] _RAND_147;
  reg [31:0] _RAND_148;
  reg [31:0] _RAND_149;
  reg [31:0] _RAND_150;
  reg [31:0] _RAND_151;
  reg [31:0] _RAND_152;
  reg [31:0] _RAND_153;
  reg [31:0] _RAND_154;
  reg [31:0] _RAND_155;
  reg [31:0] _RAND_156;
  reg [31:0] _RAND_157;
  reg [31:0] _RAND_158;
  reg [31:0] _RAND_159;
  reg [31:0] _RAND_160;
  reg [31:0] _RAND_161;
  reg [31:0] _RAND_162;
  reg [31:0] _RAND_163;
  reg [31:0] _RAND_164;
  reg [31:0] _RAND_165;
  reg [31:0] _RAND_166;
  reg [31:0] _RAND_167;
  reg [31:0] _RAND_168;
  reg [31:0] _RAND_169;
  reg [31:0] _RAND_170;
  reg [31:0] _RAND_171;
  reg [31:0] _RAND_172;
  reg [31:0] _RAND_173;
  reg [31:0] _RAND_174;
  reg [31:0] _RAND_175;
  reg [31:0] _RAND_176;
  reg [31:0] _RAND_177;
  reg [31:0] _RAND_178;
  reg [31:0] _RAND_179;
  reg [31:0] _RAND_180;
  reg [31:0] _RAND_181;
  reg [31:0] _RAND_182;
  reg [31:0] _RAND_183;
  reg [31:0] _RAND_184;
  reg [31:0] _RAND_185;
  reg [31:0] _RAND_186;
  reg [31:0] _RAND_187;
  reg [31:0] _RAND_188;
  reg [31:0] _RAND_189;
  reg [31:0] _RAND_190;
  reg [31:0] _RAND_191;
  reg [31:0] _RAND_192;
  reg [31:0] _RAND_193;
  reg [31:0] _RAND_194;
  reg [31:0] _RAND_195;
  reg [31:0] _RAND_196;
  reg [31:0] _RAND_197;
  reg [31:0] _RAND_198;
  reg [31:0] _RAND_199;
  reg [31:0] _RAND_200;
  reg [31:0] _RAND_201;
  reg [31:0] _RAND_202;
  reg [31:0] _RAND_203;
  reg [31:0] _RAND_204;
  reg [31:0] _RAND_205;
  reg [31:0] _RAND_206;
  reg [31:0] _RAND_207;
  reg [31:0] _RAND_208;
  reg [31:0] _RAND_209;
  reg [31:0] _RAND_210;
  reg [31:0] _RAND_211;
  reg [31:0] _RAND_212;
  reg [31:0] _RAND_213;
  reg [31:0] _RAND_214;
  reg [31:0] _RAND_215;
  reg [31:0] _RAND_216;
  reg [31:0] _RAND_217;
  reg [31:0] _RAND_218;
  reg [31:0] _RAND_219;
  reg [31:0] _RAND_220;
  reg [31:0] _RAND_221;
  reg [31:0] _RAND_222;
  reg [31:0] _RAND_223;
  reg [31:0] _RAND_224;
  reg [31:0] _RAND_225;
  reg [31:0] _RAND_226;
  reg [31:0] _RAND_227;
  reg [31:0] _RAND_228;
  reg [31:0] _RAND_229;
  reg [31:0] _RAND_230;
  reg [31:0] _RAND_231;
  reg [31:0] _RAND_232;
  reg [31:0] _RAND_233;
  reg [31:0] _RAND_234;
  reg [31:0] _RAND_235;
  reg [31:0] _RAND_236;
  reg [31:0] _RAND_237;
  reg [31:0] _RAND_238;
  reg [31:0] _RAND_239;
  reg [31:0] _RAND_240;
  reg [31:0] _RAND_241;
  reg [31:0] _RAND_242;
  reg [31:0] _RAND_243;
  reg [31:0] _RAND_244;
  reg [31:0] _RAND_245;
  reg [31:0] _RAND_246;
  reg [31:0] _RAND_247;
  reg [31:0] _RAND_248;
  reg [31:0] _RAND_249;
  reg [31:0] _RAND_250;
  reg [31:0] _RAND_251;
  reg [31:0] _RAND_252;
  reg [31:0] _RAND_253;
  reg [31:0] _RAND_254;
  reg [31:0] _RAND_255;
  reg [31:0] _RAND_256;
  reg [31:0] _RAND_257;
  reg [31:0] _RAND_258;
  reg [31:0] _RAND_259;
  reg [31:0] _RAND_260;
  reg [31:0] _RAND_261;
  reg [31:0] _RAND_262;
  reg [31:0] _RAND_263;
  reg [31:0] _RAND_264;
  reg [31:0] _RAND_265;
  reg [31:0] _RAND_266;
  reg [31:0] _RAND_267;
  reg [31:0] _RAND_268;
  reg [31:0] _RAND_269;
  reg [31:0] _RAND_270;
  reg [31:0] _RAND_271;
  reg [31:0] _RAND_272;
  reg [31:0] _RAND_273;
  reg [31:0] _RAND_274;
  reg [31:0] _RAND_275;
  reg [31:0] _RAND_276;
  reg [31:0] _RAND_277;
  reg [31:0] _RAND_278;
  reg [31:0] _RAND_279;
  reg [31:0] _RAND_280;
  reg [31:0] _RAND_281;
  reg [31:0] _RAND_282;
  reg [31:0] _RAND_283;
  reg [31:0] _RAND_284;
  reg [31:0] _RAND_285;
  reg [31:0] _RAND_286;
  reg [31:0] _RAND_287;
  reg [31:0] _RAND_288;
  reg [31:0] _RAND_289;
  reg [31:0] _RAND_290;
  reg [31:0] _RAND_291;
  reg [31:0] _RAND_292;
  reg [31:0] _RAND_293;
  reg [31:0] _RAND_294;
  reg [31:0] _RAND_295;
  reg [31:0] _RAND_296;
  reg [31:0] _RAND_297;
  reg [31:0] _RAND_298;
  reg [31:0] _RAND_299;
  reg [31:0] _RAND_300;
  reg [31:0] _RAND_301;
  reg [31:0] _RAND_302;
  reg [31:0] _RAND_303;
  reg [31:0] _RAND_304;
  reg [31:0] _RAND_305;
  reg [31:0] _RAND_306;
  reg [31:0] _RAND_307;
  reg [31:0] _RAND_308;
  reg [31:0] _RAND_309;
  reg [31:0] _RAND_310;
  reg [31:0] _RAND_311;
  reg [31:0] _RAND_312;
  reg [31:0] _RAND_313;
  reg [31:0] _RAND_314;
  reg [31:0] _RAND_315;
  reg [31:0] _RAND_316;
  reg [31:0] _RAND_317;
  reg [31:0] _RAND_318;
  reg [31:0] _RAND_319;
  reg [31:0] _RAND_320;
  reg [31:0] _RAND_321;
  reg [31:0] _RAND_322;
  reg [31:0] _RAND_323;
  reg [31:0] _RAND_324;
  reg [31:0] _RAND_325;
  reg [31:0] _RAND_326;
  reg [31:0] _RAND_327;
  reg [31:0] _RAND_328;
  reg [31:0] _RAND_329;
  reg [31:0] _RAND_330;
  reg [31:0] _RAND_331;
  reg [31:0] _RAND_332;
  reg [31:0] _RAND_333;
  reg [31:0] _RAND_334;
  reg [31:0] _RAND_335;
  reg [31:0] _RAND_336;
  reg [31:0] _RAND_337;
  reg [31:0] _RAND_338;
  reg [31:0] _RAND_339;
  reg [31:0] _RAND_340;
  reg [31:0] _RAND_341;
  reg [31:0] _RAND_342;
  reg [31:0] _RAND_343;
  reg [31:0] _RAND_344;
  reg [31:0] _RAND_345;
  reg [31:0] _RAND_346;
  reg [31:0] _RAND_347;
  reg [31:0] _RAND_348;
  reg [31:0] _RAND_349;
  reg [31:0] _RAND_350;
  reg [31:0] _RAND_351;
  reg [31:0] _RAND_352;
  reg [31:0] _RAND_353;
  reg [31:0] _RAND_354;
  reg [31:0] _RAND_355;
  reg [31:0] _RAND_356;
  reg [31:0] _RAND_357;
  reg [31:0] _RAND_358;
  reg [31:0] _RAND_359;
  reg [31:0] _RAND_360;
  reg [31:0] _RAND_361;
  reg [31:0] _RAND_362;
  reg [31:0] _RAND_363;
  reg [31:0] _RAND_364;
  reg [31:0] _RAND_365;
  reg [31:0] _RAND_366;
  reg [31:0] _RAND_367;
  reg [31:0] _RAND_368;
  reg [31:0] _RAND_369;
  reg [31:0] _RAND_370;
  reg [31:0] _RAND_371;
  reg [31:0] _RAND_372;
  reg [31:0] _RAND_373;
  reg [31:0] _RAND_374;
  reg [31:0] _RAND_375;
  reg [31:0] _RAND_376;
  reg [31:0] _RAND_377;
  reg [31:0] _RAND_378;
  reg [31:0] _RAND_379;
  reg [31:0] _RAND_380;
  reg [31:0] _RAND_381;
  reg [31:0] _RAND_382;
  reg [31:0] _RAND_383;
  reg [31:0] _RAND_384;
  reg [31:0] _RAND_385;
  reg [31:0] _RAND_386;
  reg [31:0] _RAND_387;
  reg [31:0] _RAND_388;
  reg [31:0] _RAND_389;
  reg [31:0] _RAND_390;
  reg [31:0] _RAND_391;
  reg [31:0] _RAND_392;
  reg [31:0] _RAND_393;
  reg [31:0] _RAND_394;
  reg [31:0] _RAND_395;
  reg [31:0] _RAND_396;
  reg [31:0] _RAND_397;
  reg [31:0] _RAND_398;
  reg [31:0] _RAND_399;
  reg [31:0] _RAND_400;
  reg [31:0] _RAND_401;
  reg [31:0] _RAND_402;
  reg [31:0] _RAND_403;
  reg [31:0] _RAND_404;
  reg [31:0] _RAND_405;
  reg [31:0] _RAND_406;
  reg [31:0] _RAND_407;
  reg [31:0] _RAND_408;
  reg [31:0] _RAND_409;
  reg [31:0] _RAND_410;
  reg [31:0] _RAND_411;
  reg [31:0] _RAND_412;
  reg [31:0] _RAND_413;
  reg [31:0] _RAND_414;
  reg [31:0] _RAND_415;
  reg [31:0] _RAND_416;
  reg [31:0] _RAND_417;
  reg [31:0] _RAND_418;
  reg [31:0] _RAND_419;
  reg [31:0] _RAND_420;
  reg [31:0] _RAND_421;
  reg [31:0] _RAND_422;
  reg [31:0] _RAND_423;
  reg [31:0] _RAND_424;
  reg [31:0] _RAND_425;
  reg [31:0] _RAND_426;
  reg [31:0] _RAND_427;
  reg [31:0] _RAND_428;
  reg [31:0] _RAND_429;
  reg [31:0] _RAND_430;
  reg [31:0] _RAND_431;
  reg [31:0] _RAND_432;
  reg [31:0] _RAND_433;
  reg [31:0] _RAND_434;
  reg [31:0] _RAND_435;
  reg [31:0] _RAND_436;
  reg [31:0] _RAND_437;
  reg [31:0] _RAND_438;
  reg [31:0] _RAND_439;
  reg [31:0] _RAND_440;
  reg [31:0] _RAND_441;
  reg [31:0] _RAND_442;
  reg [31:0] _RAND_443;
  reg [31:0] _RAND_444;
  reg [31:0] _RAND_445;
  reg [31:0] _RAND_446;
  reg [31:0] _RAND_447;
  reg [31:0] _RAND_448;
  reg [31:0] _RAND_449;
  reg [31:0] _RAND_450;
  reg [31:0] _RAND_451;
  reg [31:0] _RAND_452;
  reg [31:0] _RAND_453;
  reg [31:0] _RAND_454;
  reg [31:0] _RAND_455;
  reg [31:0] _RAND_456;
  reg [31:0] _RAND_457;
  reg [31:0] _RAND_458;
  reg [31:0] _RAND_459;
  reg [31:0] _RAND_460;
  reg [31:0] _RAND_461;
  reg [31:0] _RAND_462;
  reg [31:0] _RAND_463;
  reg [31:0] _RAND_464;
  reg [31:0] _RAND_465;
  reg [31:0] _RAND_466;
  reg [31:0] _RAND_467;
  reg [31:0] _RAND_468;
  reg [31:0] _RAND_469;
  reg [31:0] _RAND_470;
  reg [31:0] _RAND_471;
  reg [31:0] _RAND_472;
  reg [31:0] _RAND_473;
  reg [31:0] _RAND_474;
  reg [31:0] _RAND_475;
  reg [31:0] _RAND_476;
  reg [31:0] _RAND_477;
  reg [31:0] _RAND_478;
  reg [31:0] _RAND_479;
  reg [31:0] _RAND_480;
  reg [31:0] _RAND_481;
  reg [31:0] _RAND_482;
  reg [31:0] _RAND_483;
  reg [31:0] _RAND_484;
  reg [31:0] _RAND_485;
  reg [31:0] _RAND_486;
  reg [31:0] _RAND_487;
  reg [31:0] _RAND_488;
  reg [31:0] _RAND_489;
  reg [31:0] _RAND_490;
  reg [31:0] _RAND_491;
  reg [31:0] _RAND_492;
  reg [31:0] _RAND_493;
  reg [31:0] _RAND_494;
  reg [31:0] _RAND_495;
  reg [31:0] _RAND_496;
  reg [31:0] _RAND_497;
  reg [31:0] _RAND_498;
  reg [31:0] _RAND_499;
  reg [31:0] _RAND_500;
  reg [31:0] _RAND_501;
  reg [31:0] _RAND_502;
  reg [31:0] _RAND_503;
  reg [31:0] _RAND_504;
  reg [31:0] _RAND_505;
  reg [31:0] _RAND_506;
  reg [31:0] _RAND_507;
  reg [31:0] _RAND_508;
  reg [31:0] _RAND_509;
  reg [31:0] _RAND_510;
  reg [31:0] _RAND_511;
  reg [31:0] _RAND_512;
  reg [31:0] _RAND_513;
  reg [31:0] _RAND_514;
  reg [31:0] _RAND_515;
  reg [31:0] _RAND_516;
  reg [31:0] _RAND_517;
  reg [31:0] _RAND_518;
  reg [31:0] _RAND_519;
  reg [31:0] _RAND_520;
  reg [31:0] _RAND_521;
  reg [31:0] _RAND_522;
  reg [31:0] _RAND_523;
  reg [31:0] _RAND_524;
  reg [31:0] _RAND_525;
  reg [31:0] _RAND_526;
  reg [31:0] _RAND_527;
  reg [31:0] _RAND_528;
  reg [31:0] _RAND_529;
  reg [31:0] _RAND_530;
  reg [31:0] _RAND_531;
  reg [31:0] _RAND_532;
  reg [31:0] _RAND_533;
  reg [31:0] _RAND_534;
  reg [31:0] _RAND_535;
  reg [31:0] _RAND_536;
  reg [31:0] _RAND_537;
  reg [31:0] _RAND_538;
  reg [31:0] _RAND_539;
  reg [31:0] _RAND_540;
  reg [31:0] _RAND_541;
  reg [31:0] _RAND_542;
  reg [31:0] _RAND_543;
  reg [31:0] _RAND_544;
  reg [31:0] _RAND_545;
  reg [31:0] _RAND_546;
  reg [31:0] _RAND_547;
  reg [31:0] _RAND_548;
  reg [31:0] _RAND_549;
  reg [31:0] _RAND_550;
  reg [31:0] _RAND_551;
  reg [31:0] _RAND_552;
  reg [31:0] _RAND_553;
  reg [31:0] _RAND_554;
  reg [31:0] _RAND_555;
  reg [31:0] _RAND_556;
  reg [31:0] _RAND_557;
  reg [31:0] _RAND_558;
  reg [31:0] _RAND_559;
  reg [31:0] _RAND_560;
  reg [31:0] _RAND_561;
  reg [31:0] _RAND_562;
  reg [31:0] _RAND_563;
  reg [31:0] _RAND_564;
  reg [31:0] _RAND_565;
  reg [31:0] _RAND_566;
  reg [31:0] _RAND_567;
  reg [31:0] _RAND_568;
  reg [31:0] _RAND_569;
  reg [31:0] _RAND_570;
  reg [31:0] _RAND_571;
  reg [31:0] _RAND_572;
  reg [31:0] _RAND_573;
  reg [31:0] _RAND_574;
  reg [31:0] _RAND_575;
  reg [31:0] _RAND_576;
  reg [31:0] _RAND_577;
  reg [31:0] _RAND_578;
  reg [31:0] _RAND_579;
  reg [31:0] _RAND_580;
  reg [31:0] _RAND_581;
  reg [31:0] _RAND_582;
  reg [31:0] _RAND_583;
  reg [31:0] _RAND_584;
  reg [31:0] _RAND_585;
  reg [31:0] _RAND_586;
  reg [31:0] _RAND_587;
  reg [31:0] _RAND_588;
  reg [31:0] _RAND_589;
  reg [31:0] _RAND_590;
  reg [31:0] _RAND_591;
  reg [31:0] _RAND_592;
  reg [31:0] _RAND_593;
  reg [31:0] _RAND_594;
  reg [31:0] _RAND_595;
  reg [31:0] _RAND_596;
  reg [31:0] _RAND_597;
  reg [31:0] _RAND_598;
  reg [31:0] _RAND_599;
  reg [31:0] _RAND_600;
  reg [31:0] _RAND_601;
  reg [31:0] _RAND_602;
  reg [31:0] _RAND_603;
  reg [31:0] _RAND_604;
  reg [31:0] _RAND_605;
  reg [31:0] _RAND_606;
  reg [31:0] _RAND_607;
  reg [31:0] _RAND_608;
  reg [31:0] _RAND_609;
  reg [31:0] _RAND_610;
  reg [31:0] _RAND_611;
  reg [31:0] _RAND_612;
  reg [31:0] _RAND_613;
  reg [31:0] _RAND_614;
  reg [31:0] _RAND_615;
  reg [31:0] _RAND_616;
  reg [31:0] _RAND_617;
  reg [31:0] _RAND_618;
  reg [31:0] _RAND_619;
  reg [31:0] _RAND_620;
  reg [31:0] _RAND_621;
  reg [31:0] _RAND_622;
  reg [31:0] _RAND_623;
  reg [31:0] _RAND_624;
  reg [31:0] _RAND_625;
  reg [31:0] _RAND_626;
  reg [31:0] _RAND_627;
  reg [31:0] _RAND_628;
  reg [31:0] _RAND_629;
  reg [31:0] _RAND_630;
  reg [31:0] _RAND_631;
  reg [31:0] _RAND_632;
  reg [31:0] _RAND_633;
  reg [31:0] _RAND_634;
  reg [31:0] _RAND_635;
  reg [31:0] _RAND_636;
  reg [31:0] _RAND_637;
  reg [31:0] _RAND_638;
  reg [31:0] _RAND_639;
  reg [31:0] _RAND_640;
  reg [31:0] _RAND_641;
  reg [31:0] _RAND_642;
  reg [31:0] _RAND_643;
  reg [31:0] _RAND_644;
  reg [31:0] _RAND_645;
  reg [31:0] _RAND_646;
  reg [31:0] _RAND_647;
  reg [31:0] _RAND_648;
  reg [31:0] _RAND_649;
  reg [31:0] _RAND_650;
  reg [31:0] _RAND_651;
  reg [31:0] _RAND_652;
  reg [31:0] _RAND_653;
  reg [31:0] _RAND_654;
  reg [31:0] _RAND_655;
  reg [31:0] _RAND_656;
  reg [31:0] _RAND_657;
  reg [31:0] _RAND_658;
  reg [31:0] _RAND_659;
  reg [31:0] _RAND_660;
  reg [31:0] _RAND_661;
  reg [31:0] _RAND_662;
  reg [31:0] _RAND_663;
  reg [31:0] _RAND_664;
  reg [31:0] _RAND_665;
  reg [31:0] _RAND_666;
  reg [31:0] _RAND_667;
  reg [31:0] _RAND_668;
  reg [31:0] _RAND_669;
  reg [31:0] _RAND_670;
  reg [31:0] _RAND_671;
  reg [31:0] _RAND_672;
  reg [31:0] _RAND_673;
  reg [31:0] _RAND_674;
  reg [31:0] _RAND_675;
  reg [31:0] _RAND_676;
  reg [31:0] _RAND_677;
  reg [31:0] _RAND_678;
  reg [31:0] _RAND_679;
  reg [31:0] _RAND_680;
  reg [31:0] _RAND_681;
  reg [31:0] _RAND_682;
  reg [31:0] _RAND_683;
  reg [31:0] _RAND_684;
  reg [31:0] _RAND_685;
  reg [31:0] _RAND_686;
  reg [31:0] _RAND_687;
  reg [31:0] _RAND_688;
  reg [31:0] _RAND_689;
  reg [31:0] _RAND_690;
  reg [31:0] _RAND_691;
  reg [31:0] _RAND_692;
  reg [31:0] _RAND_693;
  reg [31:0] _RAND_694;
  reg [31:0] _RAND_695;
  reg [31:0] _RAND_696;
  reg [31:0] _RAND_697;
  reg [31:0] _RAND_698;
  reg [31:0] _RAND_699;
  reg [31:0] _RAND_700;
  reg [31:0] _RAND_701;
  reg [31:0] _RAND_702;
  reg [31:0] _RAND_703;
  reg [31:0] _RAND_704;
  reg [31:0] _RAND_705;
  reg [31:0] _RAND_706;
  reg [31:0] _RAND_707;
  reg [31:0] _RAND_708;
  reg [31:0] _RAND_709;
  reg [31:0] _RAND_710;
  reg [31:0] _RAND_711;
  reg [31:0] _RAND_712;
  reg [31:0] _RAND_713;
  reg [31:0] _RAND_714;
  reg [31:0] _RAND_715;
  reg [31:0] _RAND_716;
  reg [31:0] _RAND_717;
  reg [31:0] _RAND_718;
  reg [31:0] _RAND_719;
  reg [31:0] _RAND_720;
  reg [31:0] _RAND_721;
  reg [31:0] _RAND_722;
  reg [31:0] _RAND_723;
  reg [31:0] _RAND_724;
  reg [31:0] _RAND_725;
  reg [31:0] _RAND_726;
  reg [31:0] _RAND_727;
  reg [31:0] _RAND_728;
  reg [31:0] _RAND_729;
  reg [31:0] _RAND_730;
  reg [31:0] _RAND_731;
  reg [31:0] _RAND_732;
  reg [31:0] _RAND_733;
  reg [31:0] _RAND_734;
  reg [31:0] _RAND_735;
  reg [31:0] _RAND_736;
  reg [31:0] _RAND_737;
  reg [31:0] _RAND_738;
  reg [31:0] _RAND_739;
  reg [31:0] _RAND_740;
  reg [31:0] _RAND_741;
  reg [31:0] _RAND_742;
  reg [31:0] _RAND_743;
  reg [31:0] _RAND_744;
  reg [31:0] _RAND_745;
  reg [31:0] _RAND_746;
  reg [31:0] _RAND_747;
  reg [31:0] _RAND_748;
  reg [31:0] _RAND_749;
  reg [31:0] _RAND_750;
  reg [31:0] _RAND_751;
  reg [31:0] _RAND_752;
  reg [31:0] _RAND_753;
  reg [31:0] _RAND_754;
  reg [31:0] _RAND_755;
  reg [31:0] _RAND_756;
  reg [31:0] _RAND_757;
  reg [31:0] _RAND_758;
  reg [31:0] _RAND_759;
  reg [31:0] _RAND_760;
  reg [31:0] _RAND_761;
  reg [31:0] _RAND_762;
  reg [31:0] _RAND_763;
  reg [31:0] _RAND_764;
  reg [31:0] _RAND_765;
  reg [31:0] _RAND_766;
  reg [31:0] _RAND_767;
  reg [31:0] _RAND_768;
  reg [31:0] _RAND_769;
  reg [31:0] _RAND_770;
  reg [31:0] _RAND_771;
  reg [31:0] _RAND_772;
  reg [31:0] _RAND_773;
  reg [31:0] _RAND_774;
  reg [31:0] _RAND_775;
  reg [31:0] _RAND_776;
  reg [31:0] _RAND_777;
  reg [31:0] _RAND_778;
  reg [31:0] _RAND_779;
  reg [31:0] _RAND_780;
  reg [31:0] _RAND_781;
  reg [31:0] _RAND_782;
  reg [31:0] _RAND_783;
`endif // RANDOMIZE_REG_INIT
  reg [1:0] stateReg; // @[ChiselImProc.scala 62:28]
  reg [7:0] dataReg; // @[ChiselImProc.scala 64:23]
  reg [7:0] shadowReg; // @[ChiselImProc.scala 66:25]
  reg  userReg; // @[ChiselImProc.scala 67:23]
  reg  shadowUserReg; // @[ChiselImProc.scala 68:29]
  reg  lastReg; // @[ChiselImProc.scala 69:23]
  reg  shadowLastReg; // @[ChiselImProc.scala 70:29]
  wire  _T = 2'h0 == stateReg; // @[Conditional.scala 37:30]
  wire [7:0] _GEN_1 = io_enq_valid ? io_enq_bits : dataReg; // @[ChiselImProc.scala 77:37]
  wire  _GEN_2 = io_enq_valid ? io_enq_last : lastReg; // @[ChiselImProc.scala 77:37]
  wire  _T_1 = 2'h1 == stateReg; // @[Conditional.scala 37:30]
  wire  _T_2 = ~io_enq_valid; // @[ChiselImProc.scala 84:39]
  wire  _T_3 = io_deq_ready & _T_2; // @[ChiselImProc.scala 84:36]
  wire  _T_4 = io_deq_ready & io_enq_valid; // @[ChiselImProc.scala 87:42]
  wire  _T_5 = ~io_deq_ready; // @[ChiselImProc.scala 92:29]
  wire  _T_6 = _T_5 & io_enq_valid; // @[ChiselImProc.scala 92:43]
  wire [7:0] _GEN_4 = _T_6 ? io_enq_bits : shadowReg; // @[ChiselImProc.scala 92:60]
  wire  _GEN_5 = _T_6 ? io_enq_user : shadowUserReg; // @[ChiselImProc.scala 92:60]
  wire  _GEN_6 = _T_6 ? io_enq_last : shadowLastReg; // @[ChiselImProc.scala 92:60]
  wire [7:0] _GEN_8 = _T_4 ? io_enq_bits : dataReg; // @[ChiselImProc.scala 87:59]
  wire  _GEN_10 = _T_4 ? io_enq_last : lastReg; // @[ChiselImProc.scala 87:59]
  wire [7:0] _GEN_11 = _T_4 ? shadowReg : _GEN_4; // @[ChiselImProc.scala 87:59]
  wire  _GEN_12 = _T_4 ? shadowUserReg : _GEN_5; // @[ChiselImProc.scala 87:59]
  wire  _GEN_13 = _T_4 ? shadowLastReg : _GEN_6; // @[ChiselImProc.scala 87:59]
  wire [7:0] _GEN_16 = _T_3 ? dataReg : _GEN_8; // @[ChiselImProc.scala 84:54]
  wire  _GEN_17 = _T_3 ? lastReg : _GEN_10; // @[ChiselImProc.scala 84:54]
  wire [7:0] _GEN_18 = _T_3 ? shadowReg : _GEN_11; // @[ChiselImProc.scala 84:54]
  wire  _GEN_19 = _T_3 ? shadowUserReg : _GEN_12; // @[ChiselImProc.scala 84:54]
  wire  _GEN_20 = _T_3 ? shadowLastReg : _GEN_13; // @[ChiselImProc.scala 84:54]
  wire  _T_7 = 2'h2 == stateReg; // @[Conditional.scala 37:30]
  wire [7:0] _GEN_21 = io_deq_ready ? shadowReg : dataReg; // @[ChiselImProc.scala 100:37]
  wire  _GEN_23 = io_deq_ready ? shadowLastReg : lastReg; // @[ChiselImProc.scala 100:37]
  wire  _T_8 = 2'h3 == stateReg; // @[Conditional.scala 37:30]
  wire [7:0] _GEN_26 = _T_7 ? _GEN_21 : dataReg; // @[Conditional.scala 39:67]
  wire  _GEN_28 = _T_7 ? _GEN_23 : lastReg; // @[Conditional.scala 39:67]
  wire [7:0] _GEN_32 = _T_1 ? _GEN_16 : _GEN_26; // @[Conditional.scala 39:67]
  wire  _GEN_33 = _T_1 ? _GEN_17 : _GEN_28; // @[Conditional.scala 39:67]
  wire [7:0] _GEN_34 = _T_1 ? _GEN_18 : shadowReg; // @[Conditional.scala 39:67]
  wire  _GEN_35 = _T_1 ? _GEN_19 : shadowUserReg; // @[Conditional.scala 39:67]
  wire  _GEN_36 = _T_1 ? _GEN_20 : shadowLastReg; // @[Conditional.scala 39:67]
  wire [7:0] _GEN_39 = _T ? _GEN_1 : _GEN_32; // @[Conditional.scala 40:58]
  wire  _GEN_40 = _T ? _GEN_2 : _GEN_33; // @[Conditional.scala 40:58]
  wire [7:0] _GEN_41 = _T ? shadowReg : _GEN_34; // @[Conditional.scala 40:58]
  wire  _GEN_42 = _T ? shadowUserReg : _GEN_35; // @[Conditional.scala 40:58]
  wire  _GEN_43 = _T ? shadowLastReg : _GEN_36; // @[Conditional.scala 40:58]
  wire  _T_9 = stateReg == 2'h0; // @[ChiselImProc.scala 116:35]
  wire  _T_10 = stateReg == 2'h1; // @[ChiselImProc.scala 116:57]
  wire  _T_11 = _T_9 | _T_10; // @[ChiselImProc.scala 116:45]
  wire  _T_12 = stateReg == 2'h3; // @[ChiselImProc.scala 116:77]
  wire  _T_15 = stateReg == 2'h2; // @[ChiselImProc.scala 117:55]
  wire  _T_16 = _T_10 | _T_15; // @[ChiselImProc.scala 117:43]
  reg [7:0] lineBuffer_0; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_1; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_2; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_3; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_4; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_5; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_6; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_7; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_8; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_9; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_10; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_11; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_12; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_13; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_14; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_15; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_16; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_17; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_18; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_19; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_20; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_21; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_22; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_23; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_24; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_25; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_26; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_27; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_28; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_29; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_30; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_31; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_32; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_33; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_34; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_35; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_36; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_37; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_38; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_39; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_40; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_41; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_42; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_43; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_44; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_45; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_46; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_47; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_48; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_49; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_50; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_51; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_52; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_53; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_54; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_55; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_56; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_57; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_58; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_59; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_60; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_61; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_62; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_63; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_64; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_65; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_66; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_67; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_68; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_69; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_70; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_71; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_72; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_73; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_74; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_75; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_76; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_77; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_78; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_79; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_80; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_81; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_82; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_83; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_84; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_85; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_86; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_87; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_88; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_89; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_90; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_91; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_92; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_93; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_94; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_95; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_96; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_97; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_98; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_99; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_100; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_101; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_102; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_103; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_104; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_105; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_106; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_107; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_108; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_109; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_110; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_111; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_112; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_113; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_114; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_115; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_116; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_117; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_118; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_119; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_120; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_121; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_122; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_123; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_124; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_125; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_126; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_127; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_128; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_129; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_130; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_131; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_132; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_133; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_134; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_135; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_136; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_137; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_138; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_139; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_140; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_141; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_142; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_143; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_144; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_145; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_146; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_147; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_148; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_149; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_150; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_151; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_152; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_153; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_154; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_155; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_156; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_157; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_158; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_159; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_160; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_161; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_162; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_163; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_164; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_165; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_166; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_167; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_168; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_169; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_170; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_171; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_172; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_173; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_174; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_175; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_176; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_177; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_178; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_179; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_180; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_181; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_182; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_183; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_184; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_185; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_186; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_187; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_188; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_189; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_190; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_191; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_192; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_193; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_194; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_195; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_196; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_197; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_198; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_199; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_200; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_201; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_202; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_203; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_204; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_205; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_206; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_207; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_208; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_209; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_210; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_211; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_212; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_213; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_214; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_215; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_216; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_217; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_218; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_219; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_220; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_221; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_222; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_223; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_224; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_225; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_226; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_227; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_228; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_229; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_230; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_231; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_232; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_233; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_234; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_235; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_236; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_237; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_238; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_239; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_240; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_241; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_242; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_243; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_244; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_245; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_246; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_247; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_248; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_249; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_250; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_251; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_252; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_253; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_254; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_255; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_256; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_257; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_258; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_259; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_260; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_261; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_262; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_263; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_264; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_265; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_266; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_267; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_268; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_269; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_270; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_271; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_272; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_273; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_274; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_275; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_276; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_277; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_278; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_279; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_280; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_281; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_282; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_283; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_284; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_285; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_286; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_287; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_288; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_289; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_290; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_291; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_292; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_293; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_294; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_295; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_296; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_297; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_298; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_299; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_300; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_301; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_302; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_303; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_304; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_305; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_306; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_307; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_308; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_309; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_310; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_311; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_312; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_313; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_314; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_315; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_316; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_317; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_318; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_319; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_320; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_321; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_322; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_323; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_324; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_325; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_326; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_327; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_328; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_329; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_330; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_331; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_332; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_333; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_334; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_335; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_336; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_337; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_338; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_339; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_340; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_341; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_342; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_343; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_344; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_345; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_346; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_347; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_348; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_349; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_350; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_351; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_352; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_353; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_354; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_355; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_356; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_357; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_358; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_359; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_360; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_361; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_362; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_363; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_364; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_365; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_366; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_367; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_368; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_369; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_370; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_371; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_372; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_373; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_374; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_375; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_376; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_377; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_378; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_379; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_380; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_381; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_382; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_383; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_384; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_385; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_386; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_387; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_388; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_389; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_390; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_391; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_392; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_393; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_394; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_395; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_396; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_397; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_398; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_399; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_400; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_401; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_402; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_403; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_404; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_405; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_406; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_407; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_408; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_409; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_410; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_411; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_412; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_413; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_414; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_415; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_416; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_417; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_418; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_419; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_420; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_421; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_422; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_423; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_424; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_425; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_426; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_427; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_428; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_429; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_430; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_431; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_432; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_433; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_434; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_435; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_436; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_437; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_438; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_439; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_440; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_441; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_442; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_443; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_444; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_445; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_446; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_447; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_448; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_449; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_450; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_451; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_452; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_453; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_454; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_455; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_456; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_457; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_458; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_459; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_460; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_461; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_462; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_463; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_464; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_465; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_466; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_467; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_468; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_469; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_470; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_471; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_472; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_473; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_474; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_475; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_476; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_477; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_478; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_479; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_480; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_481; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_482; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_483; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_484; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_485; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_486; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_487; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_488; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_489; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_490; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_491; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_492; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_493; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_494; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_495; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_496; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_497; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_498; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_499; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_500; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_501; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_502; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_503; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_504; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_505; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_506; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_507; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_508; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_509; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_510; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_511; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_512; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_513; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_514; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_515; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_516; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_517; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_518; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_519; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_520; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_521; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_522; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_523; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_524; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_525; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_526; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_527; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_528; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_529; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_530; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_531; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_532; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_533; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_534; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_535; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_536; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_537; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_538; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_539; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_540; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_541; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_542; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_543; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_544; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_545; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_546; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_547; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_548; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_549; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_550; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_551; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_552; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_553; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_554; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_555; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_556; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_557; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_558; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_559; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_560; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_561; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_562; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_563; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_564; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_565; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_566; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_567; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_568; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_569; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_570; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_571; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_572; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_573; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_574; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_575; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_576; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_577; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_578; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_579; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_580; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_581; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_582; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_583; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_584; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_585; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_586; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_587; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_588; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_589; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_590; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_591; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_592; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_593; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_594; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_595; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_596; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_597; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_598; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_599; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_600; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_601; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_602; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_603; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_604; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_605; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_606; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_607; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_608; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_609; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_610; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_611; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_612; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_613; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_614; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_615; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_616; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_617; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_618; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_619; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_620; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_621; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_622; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_623; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_624; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_625; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_626; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_627; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_628; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_629; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_630; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_631; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_632; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_633; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_634; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_635; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_636; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_637; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_638; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_639; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_640; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_641; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_642; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_643; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_644; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_645; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_646; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_647; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_648; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_649; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_650; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_651; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_652; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_653; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_654; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_655; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_656; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_657; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_658; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_659; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_660; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_661; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_662; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_663; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_664; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_665; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_666; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_667; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_668; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_669; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_670; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_671; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_672; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_673; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_674; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_675; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_676; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_677; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_678; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_679; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_680; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_681; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_682; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_683; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_684; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_685; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_686; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_687; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_688; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_689; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_690; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_691; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_692; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_693; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_694; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_695; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_696; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_697; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_698; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_699; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_700; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_701; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_702; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_703; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_704; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_705; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_706; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_707; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_708; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_709; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_710; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_711; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_712; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_713; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_714; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_715; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_716; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_717; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_718; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_719; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_720; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_721; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_722; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_723; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_724; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_725; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_726; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_727; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_728; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_729; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_730; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_731; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_732; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_733; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_734; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_735; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_736; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_737; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_738; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_739; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_740; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_741; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_742; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_743; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_744; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_745; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_746; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_747; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_748; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_749; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_750; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_751; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_752; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_753; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_754; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_755; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_756; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_757; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_758; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_759; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_760; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_761; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_762; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_763; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_764; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_765; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_766; // @[ChiselImProc.scala 461:25]
  reg [7:0] lineBuffer_767; // @[ChiselImProc.scala 461:25]
  reg [7:0] windowBuffer_0; // @[ChiselImProc.scala 462:27]
  reg [7:0] windowBuffer_1; // @[ChiselImProc.scala 462:27]
  reg [7:0] windowBuffer_2; // @[ChiselImProc.scala 462:27]
  reg [7:0] windowBuffer_3; // @[ChiselImProc.scala 462:27]
  reg [7:0] windowBuffer_4; // @[ChiselImProc.scala 462:27]
  reg [7:0] windowBuffer_5; // @[ChiselImProc.scala 462:27]
  reg [7:0] windowBuffer_6; // @[ChiselImProc.scala 462:27]
  reg [7:0] windowBuffer_7; // @[ChiselImProc.scala 462:27]
  reg [7:0] windowBuffer_8; // @[ChiselImProc.scala 462:27]
  wire  sel = _T_16 & io_deq_ready; // @[ChiselImProc.scala 467:45]
  wire  _T_815 = windowBuffer_4 != 8'h0; // @[ChiselImProc.scala 482:43]
  wire  _T_817 = windowBuffer_0 != 8'hff; // @[ChiselImProc.scala 486:54]
  wire  _T_819 = windowBuffer_1 != 8'hff; // @[ChiselImProc.scala 486:54]
  wire  _T_820 = _T_817 & _T_819; // @[ChiselImProc.scala 486:34]
  wire  _T_821 = windowBuffer_2 != 8'hff; // @[ChiselImProc.scala 486:54]
  wire  _T_822 = _T_820 & _T_821; // @[ChiselImProc.scala 486:34]
  wire  _T_823 = windowBuffer_3 != 8'hff; // @[ChiselImProc.scala 486:54]
  wire  _T_824 = _T_822 & _T_823; // @[ChiselImProc.scala 486:34]
  wire  _T_825 = windowBuffer_4 != 8'hff; // @[ChiselImProc.scala 486:54]
  wire  _T_826 = _T_824 & _T_825; // @[ChiselImProc.scala 486:34]
  wire  _T_827 = windowBuffer_5 != 8'hff; // @[ChiselImProc.scala 486:54]
  wire  _T_828 = _T_826 & _T_827; // @[ChiselImProc.scala 486:34]
  wire  _T_829 = windowBuffer_6 != 8'hff; // @[ChiselImProc.scala 486:54]
  wire  _T_830 = _T_828 & _T_829; // @[ChiselImProc.scala 486:34]
  wire  _T_831 = windowBuffer_7 != 8'hff; // @[ChiselImProc.scala 486:54]
  wire  _T_832 = _T_830 & _T_831; // @[ChiselImProc.scala 486:34]
  wire [7:0] _T_833 = _T_832 ? 8'h0 : 8'hff; // @[ChiselImProc.scala 488:25]
  assign io_enq_ready = _T_11 | _T_12; // @[ChiselImProc.scala 116:22 ChiselImProc.scala 116:22]
  assign io_deq_valid = _T_10 | _T_15; // @[ChiselImProc.scala 117:22 ChiselImProc.scala 117:22]
  assign io_deq_bits = _T_815 ? _T_833 : 8'h0; // @[ChiselImProc.scala 492:17]
  assign io_deq_user = userReg; // @[ChiselImProc.scala 144:17 ChiselImProc.scala 114:21 ChiselImProc.scala 114:21]
  assign io_deq_last = lastReg; // @[ChiselImProc.scala 143:17 ChiselImProc.scala 113:21 ChiselImProc.scala 113:21]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  stateReg = _RAND_0[1:0];
  _RAND_1 = {1{`RANDOM}};
  dataReg = _RAND_1[7:0];
  _RAND_2 = {1{`RANDOM}};
  shadowReg = _RAND_2[7:0];
  _RAND_3 = {1{`RANDOM}};
  userReg = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  shadowUserReg = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  lastReg = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  shadowLastReg = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  lineBuffer_0 = _RAND_7[7:0];
  _RAND_8 = {1{`RANDOM}};
  lineBuffer_1 = _RAND_8[7:0];
  _RAND_9 = {1{`RANDOM}};
  lineBuffer_2 = _RAND_9[7:0];
  _RAND_10 = {1{`RANDOM}};
  lineBuffer_3 = _RAND_10[7:0];
  _RAND_11 = {1{`RANDOM}};
  lineBuffer_4 = _RAND_11[7:0];
  _RAND_12 = {1{`RANDOM}};
  lineBuffer_5 = _RAND_12[7:0];
  _RAND_13 = {1{`RANDOM}};
  lineBuffer_6 = _RAND_13[7:0];
  _RAND_14 = {1{`RANDOM}};
  lineBuffer_7 = _RAND_14[7:0];
  _RAND_15 = {1{`RANDOM}};
  lineBuffer_8 = _RAND_15[7:0];
  _RAND_16 = {1{`RANDOM}};
  lineBuffer_9 = _RAND_16[7:0];
  _RAND_17 = {1{`RANDOM}};
  lineBuffer_10 = _RAND_17[7:0];
  _RAND_18 = {1{`RANDOM}};
  lineBuffer_11 = _RAND_18[7:0];
  _RAND_19 = {1{`RANDOM}};
  lineBuffer_12 = _RAND_19[7:0];
  _RAND_20 = {1{`RANDOM}};
  lineBuffer_13 = _RAND_20[7:0];
  _RAND_21 = {1{`RANDOM}};
  lineBuffer_14 = _RAND_21[7:0];
  _RAND_22 = {1{`RANDOM}};
  lineBuffer_15 = _RAND_22[7:0];
  _RAND_23 = {1{`RANDOM}};
  lineBuffer_16 = _RAND_23[7:0];
  _RAND_24 = {1{`RANDOM}};
  lineBuffer_17 = _RAND_24[7:0];
  _RAND_25 = {1{`RANDOM}};
  lineBuffer_18 = _RAND_25[7:0];
  _RAND_26 = {1{`RANDOM}};
  lineBuffer_19 = _RAND_26[7:0];
  _RAND_27 = {1{`RANDOM}};
  lineBuffer_20 = _RAND_27[7:0];
  _RAND_28 = {1{`RANDOM}};
  lineBuffer_21 = _RAND_28[7:0];
  _RAND_29 = {1{`RANDOM}};
  lineBuffer_22 = _RAND_29[7:0];
  _RAND_30 = {1{`RANDOM}};
  lineBuffer_23 = _RAND_30[7:0];
  _RAND_31 = {1{`RANDOM}};
  lineBuffer_24 = _RAND_31[7:0];
  _RAND_32 = {1{`RANDOM}};
  lineBuffer_25 = _RAND_32[7:0];
  _RAND_33 = {1{`RANDOM}};
  lineBuffer_26 = _RAND_33[7:0];
  _RAND_34 = {1{`RANDOM}};
  lineBuffer_27 = _RAND_34[7:0];
  _RAND_35 = {1{`RANDOM}};
  lineBuffer_28 = _RAND_35[7:0];
  _RAND_36 = {1{`RANDOM}};
  lineBuffer_29 = _RAND_36[7:0];
  _RAND_37 = {1{`RANDOM}};
  lineBuffer_30 = _RAND_37[7:0];
  _RAND_38 = {1{`RANDOM}};
  lineBuffer_31 = _RAND_38[7:0];
  _RAND_39 = {1{`RANDOM}};
  lineBuffer_32 = _RAND_39[7:0];
  _RAND_40 = {1{`RANDOM}};
  lineBuffer_33 = _RAND_40[7:0];
  _RAND_41 = {1{`RANDOM}};
  lineBuffer_34 = _RAND_41[7:0];
  _RAND_42 = {1{`RANDOM}};
  lineBuffer_35 = _RAND_42[7:0];
  _RAND_43 = {1{`RANDOM}};
  lineBuffer_36 = _RAND_43[7:0];
  _RAND_44 = {1{`RANDOM}};
  lineBuffer_37 = _RAND_44[7:0];
  _RAND_45 = {1{`RANDOM}};
  lineBuffer_38 = _RAND_45[7:0];
  _RAND_46 = {1{`RANDOM}};
  lineBuffer_39 = _RAND_46[7:0];
  _RAND_47 = {1{`RANDOM}};
  lineBuffer_40 = _RAND_47[7:0];
  _RAND_48 = {1{`RANDOM}};
  lineBuffer_41 = _RAND_48[7:0];
  _RAND_49 = {1{`RANDOM}};
  lineBuffer_42 = _RAND_49[7:0];
  _RAND_50 = {1{`RANDOM}};
  lineBuffer_43 = _RAND_50[7:0];
  _RAND_51 = {1{`RANDOM}};
  lineBuffer_44 = _RAND_51[7:0];
  _RAND_52 = {1{`RANDOM}};
  lineBuffer_45 = _RAND_52[7:0];
  _RAND_53 = {1{`RANDOM}};
  lineBuffer_46 = _RAND_53[7:0];
  _RAND_54 = {1{`RANDOM}};
  lineBuffer_47 = _RAND_54[7:0];
  _RAND_55 = {1{`RANDOM}};
  lineBuffer_48 = _RAND_55[7:0];
  _RAND_56 = {1{`RANDOM}};
  lineBuffer_49 = _RAND_56[7:0];
  _RAND_57 = {1{`RANDOM}};
  lineBuffer_50 = _RAND_57[7:0];
  _RAND_58 = {1{`RANDOM}};
  lineBuffer_51 = _RAND_58[7:0];
  _RAND_59 = {1{`RANDOM}};
  lineBuffer_52 = _RAND_59[7:0];
  _RAND_60 = {1{`RANDOM}};
  lineBuffer_53 = _RAND_60[7:0];
  _RAND_61 = {1{`RANDOM}};
  lineBuffer_54 = _RAND_61[7:0];
  _RAND_62 = {1{`RANDOM}};
  lineBuffer_55 = _RAND_62[7:0];
  _RAND_63 = {1{`RANDOM}};
  lineBuffer_56 = _RAND_63[7:0];
  _RAND_64 = {1{`RANDOM}};
  lineBuffer_57 = _RAND_64[7:0];
  _RAND_65 = {1{`RANDOM}};
  lineBuffer_58 = _RAND_65[7:0];
  _RAND_66 = {1{`RANDOM}};
  lineBuffer_59 = _RAND_66[7:0];
  _RAND_67 = {1{`RANDOM}};
  lineBuffer_60 = _RAND_67[7:0];
  _RAND_68 = {1{`RANDOM}};
  lineBuffer_61 = _RAND_68[7:0];
  _RAND_69 = {1{`RANDOM}};
  lineBuffer_62 = _RAND_69[7:0];
  _RAND_70 = {1{`RANDOM}};
  lineBuffer_63 = _RAND_70[7:0];
  _RAND_71 = {1{`RANDOM}};
  lineBuffer_64 = _RAND_71[7:0];
  _RAND_72 = {1{`RANDOM}};
  lineBuffer_65 = _RAND_72[7:0];
  _RAND_73 = {1{`RANDOM}};
  lineBuffer_66 = _RAND_73[7:0];
  _RAND_74 = {1{`RANDOM}};
  lineBuffer_67 = _RAND_74[7:0];
  _RAND_75 = {1{`RANDOM}};
  lineBuffer_68 = _RAND_75[7:0];
  _RAND_76 = {1{`RANDOM}};
  lineBuffer_69 = _RAND_76[7:0];
  _RAND_77 = {1{`RANDOM}};
  lineBuffer_70 = _RAND_77[7:0];
  _RAND_78 = {1{`RANDOM}};
  lineBuffer_71 = _RAND_78[7:0];
  _RAND_79 = {1{`RANDOM}};
  lineBuffer_72 = _RAND_79[7:0];
  _RAND_80 = {1{`RANDOM}};
  lineBuffer_73 = _RAND_80[7:0];
  _RAND_81 = {1{`RANDOM}};
  lineBuffer_74 = _RAND_81[7:0];
  _RAND_82 = {1{`RANDOM}};
  lineBuffer_75 = _RAND_82[7:0];
  _RAND_83 = {1{`RANDOM}};
  lineBuffer_76 = _RAND_83[7:0];
  _RAND_84 = {1{`RANDOM}};
  lineBuffer_77 = _RAND_84[7:0];
  _RAND_85 = {1{`RANDOM}};
  lineBuffer_78 = _RAND_85[7:0];
  _RAND_86 = {1{`RANDOM}};
  lineBuffer_79 = _RAND_86[7:0];
  _RAND_87 = {1{`RANDOM}};
  lineBuffer_80 = _RAND_87[7:0];
  _RAND_88 = {1{`RANDOM}};
  lineBuffer_81 = _RAND_88[7:0];
  _RAND_89 = {1{`RANDOM}};
  lineBuffer_82 = _RAND_89[7:0];
  _RAND_90 = {1{`RANDOM}};
  lineBuffer_83 = _RAND_90[7:0];
  _RAND_91 = {1{`RANDOM}};
  lineBuffer_84 = _RAND_91[7:0];
  _RAND_92 = {1{`RANDOM}};
  lineBuffer_85 = _RAND_92[7:0];
  _RAND_93 = {1{`RANDOM}};
  lineBuffer_86 = _RAND_93[7:0];
  _RAND_94 = {1{`RANDOM}};
  lineBuffer_87 = _RAND_94[7:0];
  _RAND_95 = {1{`RANDOM}};
  lineBuffer_88 = _RAND_95[7:0];
  _RAND_96 = {1{`RANDOM}};
  lineBuffer_89 = _RAND_96[7:0];
  _RAND_97 = {1{`RANDOM}};
  lineBuffer_90 = _RAND_97[7:0];
  _RAND_98 = {1{`RANDOM}};
  lineBuffer_91 = _RAND_98[7:0];
  _RAND_99 = {1{`RANDOM}};
  lineBuffer_92 = _RAND_99[7:0];
  _RAND_100 = {1{`RANDOM}};
  lineBuffer_93 = _RAND_100[7:0];
  _RAND_101 = {1{`RANDOM}};
  lineBuffer_94 = _RAND_101[7:0];
  _RAND_102 = {1{`RANDOM}};
  lineBuffer_95 = _RAND_102[7:0];
  _RAND_103 = {1{`RANDOM}};
  lineBuffer_96 = _RAND_103[7:0];
  _RAND_104 = {1{`RANDOM}};
  lineBuffer_97 = _RAND_104[7:0];
  _RAND_105 = {1{`RANDOM}};
  lineBuffer_98 = _RAND_105[7:0];
  _RAND_106 = {1{`RANDOM}};
  lineBuffer_99 = _RAND_106[7:0];
  _RAND_107 = {1{`RANDOM}};
  lineBuffer_100 = _RAND_107[7:0];
  _RAND_108 = {1{`RANDOM}};
  lineBuffer_101 = _RAND_108[7:0];
  _RAND_109 = {1{`RANDOM}};
  lineBuffer_102 = _RAND_109[7:0];
  _RAND_110 = {1{`RANDOM}};
  lineBuffer_103 = _RAND_110[7:0];
  _RAND_111 = {1{`RANDOM}};
  lineBuffer_104 = _RAND_111[7:0];
  _RAND_112 = {1{`RANDOM}};
  lineBuffer_105 = _RAND_112[7:0];
  _RAND_113 = {1{`RANDOM}};
  lineBuffer_106 = _RAND_113[7:0];
  _RAND_114 = {1{`RANDOM}};
  lineBuffer_107 = _RAND_114[7:0];
  _RAND_115 = {1{`RANDOM}};
  lineBuffer_108 = _RAND_115[7:0];
  _RAND_116 = {1{`RANDOM}};
  lineBuffer_109 = _RAND_116[7:0];
  _RAND_117 = {1{`RANDOM}};
  lineBuffer_110 = _RAND_117[7:0];
  _RAND_118 = {1{`RANDOM}};
  lineBuffer_111 = _RAND_118[7:0];
  _RAND_119 = {1{`RANDOM}};
  lineBuffer_112 = _RAND_119[7:0];
  _RAND_120 = {1{`RANDOM}};
  lineBuffer_113 = _RAND_120[7:0];
  _RAND_121 = {1{`RANDOM}};
  lineBuffer_114 = _RAND_121[7:0];
  _RAND_122 = {1{`RANDOM}};
  lineBuffer_115 = _RAND_122[7:0];
  _RAND_123 = {1{`RANDOM}};
  lineBuffer_116 = _RAND_123[7:0];
  _RAND_124 = {1{`RANDOM}};
  lineBuffer_117 = _RAND_124[7:0];
  _RAND_125 = {1{`RANDOM}};
  lineBuffer_118 = _RAND_125[7:0];
  _RAND_126 = {1{`RANDOM}};
  lineBuffer_119 = _RAND_126[7:0];
  _RAND_127 = {1{`RANDOM}};
  lineBuffer_120 = _RAND_127[7:0];
  _RAND_128 = {1{`RANDOM}};
  lineBuffer_121 = _RAND_128[7:0];
  _RAND_129 = {1{`RANDOM}};
  lineBuffer_122 = _RAND_129[7:0];
  _RAND_130 = {1{`RANDOM}};
  lineBuffer_123 = _RAND_130[7:0];
  _RAND_131 = {1{`RANDOM}};
  lineBuffer_124 = _RAND_131[7:0];
  _RAND_132 = {1{`RANDOM}};
  lineBuffer_125 = _RAND_132[7:0];
  _RAND_133 = {1{`RANDOM}};
  lineBuffer_126 = _RAND_133[7:0];
  _RAND_134 = {1{`RANDOM}};
  lineBuffer_127 = _RAND_134[7:0];
  _RAND_135 = {1{`RANDOM}};
  lineBuffer_128 = _RAND_135[7:0];
  _RAND_136 = {1{`RANDOM}};
  lineBuffer_129 = _RAND_136[7:0];
  _RAND_137 = {1{`RANDOM}};
  lineBuffer_130 = _RAND_137[7:0];
  _RAND_138 = {1{`RANDOM}};
  lineBuffer_131 = _RAND_138[7:0];
  _RAND_139 = {1{`RANDOM}};
  lineBuffer_132 = _RAND_139[7:0];
  _RAND_140 = {1{`RANDOM}};
  lineBuffer_133 = _RAND_140[7:0];
  _RAND_141 = {1{`RANDOM}};
  lineBuffer_134 = _RAND_141[7:0];
  _RAND_142 = {1{`RANDOM}};
  lineBuffer_135 = _RAND_142[7:0];
  _RAND_143 = {1{`RANDOM}};
  lineBuffer_136 = _RAND_143[7:0];
  _RAND_144 = {1{`RANDOM}};
  lineBuffer_137 = _RAND_144[7:0];
  _RAND_145 = {1{`RANDOM}};
  lineBuffer_138 = _RAND_145[7:0];
  _RAND_146 = {1{`RANDOM}};
  lineBuffer_139 = _RAND_146[7:0];
  _RAND_147 = {1{`RANDOM}};
  lineBuffer_140 = _RAND_147[7:0];
  _RAND_148 = {1{`RANDOM}};
  lineBuffer_141 = _RAND_148[7:0];
  _RAND_149 = {1{`RANDOM}};
  lineBuffer_142 = _RAND_149[7:0];
  _RAND_150 = {1{`RANDOM}};
  lineBuffer_143 = _RAND_150[7:0];
  _RAND_151 = {1{`RANDOM}};
  lineBuffer_144 = _RAND_151[7:0];
  _RAND_152 = {1{`RANDOM}};
  lineBuffer_145 = _RAND_152[7:0];
  _RAND_153 = {1{`RANDOM}};
  lineBuffer_146 = _RAND_153[7:0];
  _RAND_154 = {1{`RANDOM}};
  lineBuffer_147 = _RAND_154[7:0];
  _RAND_155 = {1{`RANDOM}};
  lineBuffer_148 = _RAND_155[7:0];
  _RAND_156 = {1{`RANDOM}};
  lineBuffer_149 = _RAND_156[7:0];
  _RAND_157 = {1{`RANDOM}};
  lineBuffer_150 = _RAND_157[7:0];
  _RAND_158 = {1{`RANDOM}};
  lineBuffer_151 = _RAND_158[7:0];
  _RAND_159 = {1{`RANDOM}};
  lineBuffer_152 = _RAND_159[7:0];
  _RAND_160 = {1{`RANDOM}};
  lineBuffer_153 = _RAND_160[7:0];
  _RAND_161 = {1{`RANDOM}};
  lineBuffer_154 = _RAND_161[7:0];
  _RAND_162 = {1{`RANDOM}};
  lineBuffer_155 = _RAND_162[7:0];
  _RAND_163 = {1{`RANDOM}};
  lineBuffer_156 = _RAND_163[7:0];
  _RAND_164 = {1{`RANDOM}};
  lineBuffer_157 = _RAND_164[7:0];
  _RAND_165 = {1{`RANDOM}};
  lineBuffer_158 = _RAND_165[7:0];
  _RAND_166 = {1{`RANDOM}};
  lineBuffer_159 = _RAND_166[7:0];
  _RAND_167 = {1{`RANDOM}};
  lineBuffer_160 = _RAND_167[7:0];
  _RAND_168 = {1{`RANDOM}};
  lineBuffer_161 = _RAND_168[7:0];
  _RAND_169 = {1{`RANDOM}};
  lineBuffer_162 = _RAND_169[7:0];
  _RAND_170 = {1{`RANDOM}};
  lineBuffer_163 = _RAND_170[7:0];
  _RAND_171 = {1{`RANDOM}};
  lineBuffer_164 = _RAND_171[7:0];
  _RAND_172 = {1{`RANDOM}};
  lineBuffer_165 = _RAND_172[7:0];
  _RAND_173 = {1{`RANDOM}};
  lineBuffer_166 = _RAND_173[7:0];
  _RAND_174 = {1{`RANDOM}};
  lineBuffer_167 = _RAND_174[7:0];
  _RAND_175 = {1{`RANDOM}};
  lineBuffer_168 = _RAND_175[7:0];
  _RAND_176 = {1{`RANDOM}};
  lineBuffer_169 = _RAND_176[7:0];
  _RAND_177 = {1{`RANDOM}};
  lineBuffer_170 = _RAND_177[7:0];
  _RAND_178 = {1{`RANDOM}};
  lineBuffer_171 = _RAND_178[7:0];
  _RAND_179 = {1{`RANDOM}};
  lineBuffer_172 = _RAND_179[7:0];
  _RAND_180 = {1{`RANDOM}};
  lineBuffer_173 = _RAND_180[7:0];
  _RAND_181 = {1{`RANDOM}};
  lineBuffer_174 = _RAND_181[7:0];
  _RAND_182 = {1{`RANDOM}};
  lineBuffer_175 = _RAND_182[7:0];
  _RAND_183 = {1{`RANDOM}};
  lineBuffer_176 = _RAND_183[7:0];
  _RAND_184 = {1{`RANDOM}};
  lineBuffer_177 = _RAND_184[7:0];
  _RAND_185 = {1{`RANDOM}};
  lineBuffer_178 = _RAND_185[7:0];
  _RAND_186 = {1{`RANDOM}};
  lineBuffer_179 = _RAND_186[7:0];
  _RAND_187 = {1{`RANDOM}};
  lineBuffer_180 = _RAND_187[7:0];
  _RAND_188 = {1{`RANDOM}};
  lineBuffer_181 = _RAND_188[7:0];
  _RAND_189 = {1{`RANDOM}};
  lineBuffer_182 = _RAND_189[7:0];
  _RAND_190 = {1{`RANDOM}};
  lineBuffer_183 = _RAND_190[7:0];
  _RAND_191 = {1{`RANDOM}};
  lineBuffer_184 = _RAND_191[7:0];
  _RAND_192 = {1{`RANDOM}};
  lineBuffer_185 = _RAND_192[7:0];
  _RAND_193 = {1{`RANDOM}};
  lineBuffer_186 = _RAND_193[7:0];
  _RAND_194 = {1{`RANDOM}};
  lineBuffer_187 = _RAND_194[7:0];
  _RAND_195 = {1{`RANDOM}};
  lineBuffer_188 = _RAND_195[7:0];
  _RAND_196 = {1{`RANDOM}};
  lineBuffer_189 = _RAND_196[7:0];
  _RAND_197 = {1{`RANDOM}};
  lineBuffer_190 = _RAND_197[7:0];
  _RAND_198 = {1{`RANDOM}};
  lineBuffer_191 = _RAND_198[7:0];
  _RAND_199 = {1{`RANDOM}};
  lineBuffer_192 = _RAND_199[7:0];
  _RAND_200 = {1{`RANDOM}};
  lineBuffer_193 = _RAND_200[7:0];
  _RAND_201 = {1{`RANDOM}};
  lineBuffer_194 = _RAND_201[7:0];
  _RAND_202 = {1{`RANDOM}};
  lineBuffer_195 = _RAND_202[7:0];
  _RAND_203 = {1{`RANDOM}};
  lineBuffer_196 = _RAND_203[7:0];
  _RAND_204 = {1{`RANDOM}};
  lineBuffer_197 = _RAND_204[7:0];
  _RAND_205 = {1{`RANDOM}};
  lineBuffer_198 = _RAND_205[7:0];
  _RAND_206 = {1{`RANDOM}};
  lineBuffer_199 = _RAND_206[7:0];
  _RAND_207 = {1{`RANDOM}};
  lineBuffer_200 = _RAND_207[7:0];
  _RAND_208 = {1{`RANDOM}};
  lineBuffer_201 = _RAND_208[7:0];
  _RAND_209 = {1{`RANDOM}};
  lineBuffer_202 = _RAND_209[7:0];
  _RAND_210 = {1{`RANDOM}};
  lineBuffer_203 = _RAND_210[7:0];
  _RAND_211 = {1{`RANDOM}};
  lineBuffer_204 = _RAND_211[7:0];
  _RAND_212 = {1{`RANDOM}};
  lineBuffer_205 = _RAND_212[7:0];
  _RAND_213 = {1{`RANDOM}};
  lineBuffer_206 = _RAND_213[7:0];
  _RAND_214 = {1{`RANDOM}};
  lineBuffer_207 = _RAND_214[7:0];
  _RAND_215 = {1{`RANDOM}};
  lineBuffer_208 = _RAND_215[7:0];
  _RAND_216 = {1{`RANDOM}};
  lineBuffer_209 = _RAND_216[7:0];
  _RAND_217 = {1{`RANDOM}};
  lineBuffer_210 = _RAND_217[7:0];
  _RAND_218 = {1{`RANDOM}};
  lineBuffer_211 = _RAND_218[7:0];
  _RAND_219 = {1{`RANDOM}};
  lineBuffer_212 = _RAND_219[7:0];
  _RAND_220 = {1{`RANDOM}};
  lineBuffer_213 = _RAND_220[7:0];
  _RAND_221 = {1{`RANDOM}};
  lineBuffer_214 = _RAND_221[7:0];
  _RAND_222 = {1{`RANDOM}};
  lineBuffer_215 = _RAND_222[7:0];
  _RAND_223 = {1{`RANDOM}};
  lineBuffer_216 = _RAND_223[7:0];
  _RAND_224 = {1{`RANDOM}};
  lineBuffer_217 = _RAND_224[7:0];
  _RAND_225 = {1{`RANDOM}};
  lineBuffer_218 = _RAND_225[7:0];
  _RAND_226 = {1{`RANDOM}};
  lineBuffer_219 = _RAND_226[7:0];
  _RAND_227 = {1{`RANDOM}};
  lineBuffer_220 = _RAND_227[7:0];
  _RAND_228 = {1{`RANDOM}};
  lineBuffer_221 = _RAND_228[7:0];
  _RAND_229 = {1{`RANDOM}};
  lineBuffer_222 = _RAND_229[7:0];
  _RAND_230 = {1{`RANDOM}};
  lineBuffer_223 = _RAND_230[7:0];
  _RAND_231 = {1{`RANDOM}};
  lineBuffer_224 = _RAND_231[7:0];
  _RAND_232 = {1{`RANDOM}};
  lineBuffer_225 = _RAND_232[7:0];
  _RAND_233 = {1{`RANDOM}};
  lineBuffer_226 = _RAND_233[7:0];
  _RAND_234 = {1{`RANDOM}};
  lineBuffer_227 = _RAND_234[7:0];
  _RAND_235 = {1{`RANDOM}};
  lineBuffer_228 = _RAND_235[7:0];
  _RAND_236 = {1{`RANDOM}};
  lineBuffer_229 = _RAND_236[7:0];
  _RAND_237 = {1{`RANDOM}};
  lineBuffer_230 = _RAND_237[7:0];
  _RAND_238 = {1{`RANDOM}};
  lineBuffer_231 = _RAND_238[7:0];
  _RAND_239 = {1{`RANDOM}};
  lineBuffer_232 = _RAND_239[7:0];
  _RAND_240 = {1{`RANDOM}};
  lineBuffer_233 = _RAND_240[7:0];
  _RAND_241 = {1{`RANDOM}};
  lineBuffer_234 = _RAND_241[7:0];
  _RAND_242 = {1{`RANDOM}};
  lineBuffer_235 = _RAND_242[7:0];
  _RAND_243 = {1{`RANDOM}};
  lineBuffer_236 = _RAND_243[7:0];
  _RAND_244 = {1{`RANDOM}};
  lineBuffer_237 = _RAND_244[7:0];
  _RAND_245 = {1{`RANDOM}};
  lineBuffer_238 = _RAND_245[7:0];
  _RAND_246 = {1{`RANDOM}};
  lineBuffer_239 = _RAND_246[7:0];
  _RAND_247 = {1{`RANDOM}};
  lineBuffer_240 = _RAND_247[7:0];
  _RAND_248 = {1{`RANDOM}};
  lineBuffer_241 = _RAND_248[7:0];
  _RAND_249 = {1{`RANDOM}};
  lineBuffer_242 = _RAND_249[7:0];
  _RAND_250 = {1{`RANDOM}};
  lineBuffer_243 = _RAND_250[7:0];
  _RAND_251 = {1{`RANDOM}};
  lineBuffer_244 = _RAND_251[7:0];
  _RAND_252 = {1{`RANDOM}};
  lineBuffer_245 = _RAND_252[7:0];
  _RAND_253 = {1{`RANDOM}};
  lineBuffer_246 = _RAND_253[7:0];
  _RAND_254 = {1{`RANDOM}};
  lineBuffer_247 = _RAND_254[7:0];
  _RAND_255 = {1{`RANDOM}};
  lineBuffer_248 = _RAND_255[7:0];
  _RAND_256 = {1{`RANDOM}};
  lineBuffer_249 = _RAND_256[7:0];
  _RAND_257 = {1{`RANDOM}};
  lineBuffer_250 = _RAND_257[7:0];
  _RAND_258 = {1{`RANDOM}};
  lineBuffer_251 = _RAND_258[7:0];
  _RAND_259 = {1{`RANDOM}};
  lineBuffer_252 = _RAND_259[7:0];
  _RAND_260 = {1{`RANDOM}};
  lineBuffer_253 = _RAND_260[7:0];
  _RAND_261 = {1{`RANDOM}};
  lineBuffer_254 = _RAND_261[7:0];
  _RAND_262 = {1{`RANDOM}};
  lineBuffer_255 = _RAND_262[7:0];
  _RAND_263 = {1{`RANDOM}};
  lineBuffer_256 = _RAND_263[7:0];
  _RAND_264 = {1{`RANDOM}};
  lineBuffer_257 = _RAND_264[7:0];
  _RAND_265 = {1{`RANDOM}};
  lineBuffer_258 = _RAND_265[7:0];
  _RAND_266 = {1{`RANDOM}};
  lineBuffer_259 = _RAND_266[7:0];
  _RAND_267 = {1{`RANDOM}};
  lineBuffer_260 = _RAND_267[7:0];
  _RAND_268 = {1{`RANDOM}};
  lineBuffer_261 = _RAND_268[7:0];
  _RAND_269 = {1{`RANDOM}};
  lineBuffer_262 = _RAND_269[7:0];
  _RAND_270 = {1{`RANDOM}};
  lineBuffer_263 = _RAND_270[7:0];
  _RAND_271 = {1{`RANDOM}};
  lineBuffer_264 = _RAND_271[7:0];
  _RAND_272 = {1{`RANDOM}};
  lineBuffer_265 = _RAND_272[7:0];
  _RAND_273 = {1{`RANDOM}};
  lineBuffer_266 = _RAND_273[7:0];
  _RAND_274 = {1{`RANDOM}};
  lineBuffer_267 = _RAND_274[7:0];
  _RAND_275 = {1{`RANDOM}};
  lineBuffer_268 = _RAND_275[7:0];
  _RAND_276 = {1{`RANDOM}};
  lineBuffer_269 = _RAND_276[7:0];
  _RAND_277 = {1{`RANDOM}};
  lineBuffer_270 = _RAND_277[7:0];
  _RAND_278 = {1{`RANDOM}};
  lineBuffer_271 = _RAND_278[7:0];
  _RAND_279 = {1{`RANDOM}};
  lineBuffer_272 = _RAND_279[7:0];
  _RAND_280 = {1{`RANDOM}};
  lineBuffer_273 = _RAND_280[7:0];
  _RAND_281 = {1{`RANDOM}};
  lineBuffer_274 = _RAND_281[7:0];
  _RAND_282 = {1{`RANDOM}};
  lineBuffer_275 = _RAND_282[7:0];
  _RAND_283 = {1{`RANDOM}};
  lineBuffer_276 = _RAND_283[7:0];
  _RAND_284 = {1{`RANDOM}};
  lineBuffer_277 = _RAND_284[7:0];
  _RAND_285 = {1{`RANDOM}};
  lineBuffer_278 = _RAND_285[7:0];
  _RAND_286 = {1{`RANDOM}};
  lineBuffer_279 = _RAND_286[7:0];
  _RAND_287 = {1{`RANDOM}};
  lineBuffer_280 = _RAND_287[7:0];
  _RAND_288 = {1{`RANDOM}};
  lineBuffer_281 = _RAND_288[7:0];
  _RAND_289 = {1{`RANDOM}};
  lineBuffer_282 = _RAND_289[7:0];
  _RAND_290 = {1{`RANDOM}};
  lineBuffer_283 = _RAND_290[7:0];
  _RAND_291 = {1{`RANDOM}};
  lineBuffer_284 = _RAND_291[7:0];
  _RAND_292 = {1{`RANDOM}};
  lineBuffer_285 = _RAND_292[7:0];
  _RAND_293 = {1{`RANDOM}};
  lineBuffer_286 = _RAND_293[7:0];
  _RAND_294 = {1{`RANDOM}};
  lineBuffer_287 = _RAND_294[7:0];
  _RAND_295 = {1{`RANDOM}};
  lineBuffer_288 = _RAND_295[7:0];
  _RAND_296 = {1{`RANDOM}};
  lineBuffer_289 = _RAND_296[7:0];
  _RAND_297 = {1{`RANDOM}};
  lineBuffer_290 = _RAND_297[7:0];
  _RAND_298 = {1{`RANDOM}};
  lineBuffer_291 = _RAND_298[7:0];
  _RAND_299 = {1{`RANDOM}};
  lineBuffer_292 = _RAND_299[7:0];
  _RAND_300 = {1{`RANDOM}};
  lineBuffer_293 = _RAND_300[7:0];
  _RAND_301 = {1{`RANDOM}};
  lineBuffer_294 = _RAND_301[7:0];
  _RAND_302 = {1{`RANDOM}};
  lineBuffer_295 = _RAND_302[7:0];
  _RAND_303 = {1{`RANDOM}};
  lineBuffer_296 = _RAND_303[7:0];
  _RAND_304 = {1{`RANDOM}};
  lineBuffer_297 = _RAND_304[7:0];
  _RAND_305 = {1{`RANDOM}};
  lineBuffer_298 = _RAND_305[7:0];
  _RAND_306 = {1{`RANDOM}};
  lineBuffer_299 = _RAND_306[7:0];
  _RAND_307 = {1{`RANDOM}};
  lineBuffer_300 = _RAND_307[7:0];
  _RAND_308 = {1{`RANDOM}};
  lineBuffer_301 = _RAND_308[7:0];
  _RAND_309 = {1{`RANDOM}};
  lineBuffer_302 = _RAND_309[7:0];
  _RAND_310 = {1{`RANDOM}};
  lineBuffer_303 = _RAND_310[7:0];
  _RAND_311 = {1{`RANDOM}};
  lineBuffer_304 = _RAND_311[7:0];
  _RAND_312 = {1{`RANDOM}};
  lineBuffer_305 = _RAND_312[7:0];
  _RAND_313 = {1{`RANDOM}};
  lineBuffer_306 = _RAND_313[7:0];
  _RAND_314 = {1{`RANDOM}};
  lineBuffer_307 = _RAND_314[7:0];
  _RAND_315 = {1{`RANDOM}};
  lineBuffer_308 = _RAND_315[7:0];
  _RAND_316 = {1{`RANDOM}};
  lineBuffer_309 = _RAND_316[7:0];
  _RAND_317 = {1{`RANDOM}};
  lineBuffer_310 = _RAND_317[7:0];
  _RAND_318 = {1{`RANDOM}};
  lineBuffer_311 = _RAND_318[7:0];
  _RAND_319 = {1{`RANDOM}};
  lineBuffer_312 = _RAND_319[7:0];
  _RAND_320 = {1{`RANDOM}};
  lineBuffer_313 = _RAND_320[7:0];
  _RAND_321 = {1{`RANDOM}};
  lineBuffer_314 = _RAND_321[7:0];
  _RAND_322 = {1{`RANDOM}};
  lineBuffer_315 = _RAND_322[7:0];
  _RAND_323 = {1{`RANDOM}};
  lineBuffer_316 = _RAND_323[7:0];
  _RAND_324 = {1{`RANDOM}};
  lineBuffer_317 = _RAND_324[7:0];
  _RAND_325 = {1{`RANDOM}};
  lineBuffer_318 = _RAND_325[7:0];
  _RAND_326 = {1{`RANDOM}};
  lineBuffer_319 = _RAND_326[7:0];
  _RAND_327 = {1{`RANDOM}};
  lineBuffer_320 = _RAND_327[7:0];
  _RAND_328 = {1{`RANDOM}};
  lineBuffer_321 = _RAND_328[7:0];
  _RAND_329 = {1{`RANDOM}};
  lineBuffer_322 = _RAND_329[7:0];
  _RAND_330 = {1{`RANDOM}};
  lineBuffer_323 = _RAND_330[7:0];
  _RAND_331 = {1{`RANDOM}};
  lineBuffer_324 = _RAND_331[7:0];
  _RAND_332 = {1{`RANDOM}};
  lineBuffer_325 = _RAND_332[7:0];
  _RAND_333 = {1{`RANDOM}};
  lineBuffer_326 = _RAND_333[7:0];
  _RAND_334 = {1{`RANDOM}};
  lineBuffer_327 = _RAND_334[7:0];
  _RAND_335 = {1{`RANDOM}};
  lineBuffer_328 = _RAND_335[7:0];
  _RAND_336 = {1{`RANDOM}};
  lineBuffer_329 = _RAND_336[7:0];
  _RAND_337 = {1{`RANDOM}};
  lineBuffer_330 = _RAND_337[7:0];
  _RAND_338 = {1{`RANDOM}};
  lineBuffer_331 = _RAND_338[7:0];
  _RAND_339 = {1{`RANDOM}};
  lineBuffer_332 = _RAND_339[7:0];
  _RAND_340 = {1{`RANDOM}};
  lineBuffer_333 = _RAND_340[7:0];
  _RAND_341 = {1{`RANDOM}};
  lineBuffer_334 = _RAND_341[7:0];
  _RAND_342 = {1{`RANDOM}};
  lineBuffer_335 = _RAND_342[7:0];
  _RAND_343 = {1{`RANDOM}};
  lineBuffer_336 = _RAND_343[7:0];
  _RAND_344 = {1{`RANDOM}};
  lineBuffer_337 = _RAND_344[7:0];
  _RAND_345 = {1{`RANDOM}};
  lineBuffer_338 = _RAND_345[7:0];
  _RAND_346 = {1{`RANDOM}};
  lineBuffer_339 = _RAND_346[7:0];
  _RAND_347 = {1{`RANDOM}};
  lineBuffer_340 = _RAND_347[7:0];
  _RAND_348 = {1{`RANDOM}};
  lineBuffer_341 = _RAND_348[7:0];
  _RAND_349 = {1{`RANDOM}};
  lineBuffer_342 = _RAND_349[7:0];
  _RAND_350 = {1{`RANDOM}};
  lineBuffer_343 = _RAND_350[7:0];
  _RAND_351 = {1{`RANDOM}};
  lineBuffer_344 = _RAND_351[7:0];
  _RAND_352 = {1{`RANDOM}};
  lineBuffer_345 = _RAND_352[7:0];
  _RAND_353 = {1{`RANDOM}};
  lineBuffer_346 = _RAND_353[7:0];
  _RAND_354 = {1{`RANDOM}};
  lineBuffer_347 = _RAND_354[7:0];
  _RAND_355 = {1{`RANDOM}};
  lineBuffer_348 = _RAND_355[7:0];
  _RAND_356 = {1{`RANDOM}};
  lineBuffer_349 = _RAND_356[7:0];
  _RAND_357 = {1{`RANDOM}};
  lineBuffer_350 = _RAND_357[7:0];
  _RAND_358 = {1{`RANDOM}};
  lineBuffer_351 = _RAND_358[7:0];
  _RAND_359 = {1{`RANDOM}};
  lineBuffer_352 = _RAND_359[7:0];
  _RAND_360 = {1{`RANDOM}};
  lineBuffer_353 = _RAND_360[7:0];
  _RAND_361 = {1{`RANDOM}};
  lineBuffer_354 = _RAND_361[7:0];
  _RAND_362 = {1{`RANDOM}};
  lineBuffer_355 = _RAND_362[7:0];
  _RAND_363 = {1{`RANDOM}};
  lineBuffer_356 = _RAND_363[7:0];
  _RAND_364 = {1{`RANDOM}};
  lineBuffer_357 = _RAND_364[7:0];
  _RAND_365 = {1{`RANDOM}};
  lineBuffer_358 = _RAND_365[7:0];
  _RAND_366 = {1{`RANDOM}};
  lineBuffer_359 = _RAND_366[7:0];
  _RAND_367 = {1{`RANDOM}};
  lineBuffer_360 = _RAND_367[7:0];
  _RAND_368 = {1{`RANDOM}};
  lineBuffer_361 = _RAND_368[7:0];
  _RAND_369 = {1{`RANDOM}};
  lineBuffer_362 = _RAND_369[7:0];
  _RAND_370 = {1{`RANDOM}};
  lineBuffer_363 = _RAND_370[7:0];
  _RAND_371 = {1{`RANDOM}};
  lineBuffer_364 = _RAND_371[7:0];
  _RAND_372 = {1{`RANDOM}};
  lineBuffer_365 = _RAND_372[7:0];
  _RAND_373 = {1{`RANDOM}};
  lineBuffer_366 = _RAND_373[7:0];
  _RAND_374 = {1{`RANDOM}};
  lineBuffer_367 = _RAND_374[7:0];
  _RAND_375 = {1{`RANDOM}};
  lineBuffer_368 = _RAND_375[7:0];
  _RAND_376 = {1{`RANDOM}};
  lineBuffer_369 = _RAND_376[7:0];
  _RAND_377 = {1{`RANDOM}};
  lineBuffer_370 = _RAND_377[7:0];
  _RAND_378 = {1{`RANDOM}};
  lineBuffer_371 = _RAND_378[7:0];
  _RAND_379 = {1{`RANDOM}};
  lineBuffer_372 = _RAND_379[7:0];
  _RAND_380 = {1{`RANDOM}};
  lineBuffer_373 = _RAND_380[7:0];
  _RAND_381 = {1{`RANDOM}};
  lineBuffer_374 = _RAND_381[7:0];
  _RAND_382 = {1{`RANDOM}};
  lineBuffer_375 = _RAND_382[7:0];
  _RAND_383 = {1{`RANDOM}};
  lineBuffer_376 = _RAND_383[7:0];
  _RAND_384 = {1{`RANDOM}};
  lineBuffer_377 = _RAND_384[7:0];
  _RAND_385 = {1{`RANDOM}};
  lineBuffer_378 = _RAND_385[7:0];
  _RAND_386 = {1{`RANDOM}};
  lineBuffer_379 = _RAND_386[7:0];
  _RAND_387 = {1{`RANDOM}};
  lineBuffer_380 = _RAND_387[7:0];
  _RAND_388 = {1{`RANDOM}};
  lineBuffer_381 = _RAND_388[7:0];
  _RAND_389 = {1{`RANDOM}};
  lineBuffer_382 = _RAND_389[7:0];
  _RAND_390 = {1{`RANDOM}};
  lineBuffer_383 = _RAND_390[7:0];
  _RAND_391 = {1{`RANDOM}};
  lineBuffer_384 = _RAND_391[7:0];
  _RAND_392 = {1{`RANDOM}};
  lineBuffer_385 = _RAND_392[7:0];
  _RAND_393 = {1{`RANDOM}};
  lineBuffer_386 = _RAND_393[7:0];
  _RAND_394 = {1{`RANDOM}};
  lineBuffer_387 = _RAND_394[7:0];
  _RAND_395 = {1{`RANDOM}};
  lineBuffer_388 = _RAND_395[7:0];
  _RAND_396 = {1{`RANDOM}};
  lineBuffer_389 = _RAND_396[7:0];
  _RAND_397 = {1{`RANDOM}};
  lineBuffer_390 = _RAND_397[7:0];
  _RAND_398 = {1{`RANDOM}};
  lineBuffer_391 = _RAND_398[7:0];
  _RAND_399 = {1{`RANDOM}};
  lineBuffer_392 = _RAND_399[7:0];
  _RAND_400 = {1{`RANDOM}};
  lineBuffer_393 = _RAND_400[7:0];
  _RAND_401 = {1{`RANDOM}};
  lineBuffer_394 = _RAND_401[7:0];
  _RAND_402 = {1{`RANDOM}};
  lineBuffer_395 = _RAND_402[7:0];
  _RAND_403 = {1{`RANDOM}};
  lineBuffer_396 = _RAND_403[7:0];
  _RAND_404 = {1{`RANDOM}};
  lineBuffer_397 = _RAND_404[7:0];
  _RAND_405 = {1{`RANDOM}};
  lineBuffer_398 = _RAND_405[7:0];
  _RAND_406 = {1{`RANDOM}};
  lineBuffer_399 = _RAND_406[7:0];
  _RAND_407 = {1{`RANDOM}};
  lineBuffer_400 = _RAND_407[7:0];
  _RAND_408 = {1{`RANDOM}};
  lineBuffer_401 = _RAND_408[7:0];
  _RAND_409 = {1{`RANDOM}};
  lineBuffer_402 = _RAND_409[7:0];
  _RAND_410 = {1{`RANDOM}};
  lineBuffer_403 = _RAND_410[7:0];
  _RAND_411 = {1{`RANDOM}};
  lineBuffer_404 = _RAND_411[7:0];
  _RAND_412 = {1{`RANDOM}};
  lineBuffer_405 = _RAND_412[7:0];
  _RAND_413 = {1{`RANDOM}};
  lineBuffer_406 = _RAND_413[7:0];
  _RAND_414 = {1{`RANDOM}};
  lineBuffer_407 = _RAND_414[7:0];
  _RAND_415 = {1{`RANDOM}};
  lineBuffer_408 = _RAND_415[7:0];
  _RAND_416 = {1{`RANDOM}};
  lineBuffer_409 = _RAND_416[7:0];
  _RAND_417 = {1{`RANDOM}};
  lineBuffer_410 = _RAND_417[7:0];
  _RAND_418 = {1{`RANDOM}};
  lineBuffer_411 = _RAND_418[7:0];
  _RAND_419 = {1{`RANDOM}};
  lineBuffer_412 = _RAND_419[7:0];
  _RAND_420 = {1{`RANDOM}};
  lineBuffer_413 = _RAND_420[7:0];
  _RAND_421 = {1{`RANDOM}};
  lineBuffer_414 = _RAND_421[7:0];
  _RAND_422 = {1{`RANDOM}};
  lineBuffer_415 = _RAND_422[7:0];
  _RAND_423 = {1{`RANDOM}};
  lineBuffer_416 = _RAND_423[7:0];
  _RAND_424 = {1{`RANDOM}};
  lineBuffer_417 = _RAND_424[7:0];
  _RAND_425 = {1{`RANDOM}};
  lineBuffer_418 = _RAND_425[7:0];
  _RAND_426 = {1{`RANDOM}};
  lineBuffer_419 = _RAND_426[7:0];
  _RAND_427 = {1{`RANDOM}};
  lineBuffer_420 = _RAND_427[7:0];
  _RAND_428 = {1{`RANDOM}};
  lineBuffer_421 = _RAND_428[7:0];
  _RAND_429 = {1{`RANDOM}};
  lineBuffer_422 = _RAND_429[7:0];
  _RAND_430 = {1{`RANDOM}};
  lineBuffer_423 = _RAND_430[7:0];
  _RAND_431 = {1{`RANDOM}};
  lineBuffer_424 = _RAND_431[7:0];
  _RAND_432 = {1{`RANDOM}};
  lineBuffer_425 = _RAND_432[7:0];
  _RAND_433 = {1{`RANDOM}};
  lineBuffer_426 = _RAND_433[7:0];
  _RAND_434 = {1{`RANDOM}};
  lineBuffer_427 = _RAND_434[7:0];
  _RAND_435 = {1{`RANDOM}};
  lineBuffer_428 = _RAND_435[7:0];
  _RAND_436 = {1{`RANDOM}};
  lineBuffer_429 = _RAND_436[7:0];
  _RAND_437 = {1{`RANDOM}};
  lineBuffer_430 = _RAND_437[7:0];
  _RAND_438 = {1{`RANDOM}};
  lineBuffer_431 = _RAND_438[7:0];
  _RAND_439 = {1{`RANDOM}};
  lineBuffer_432 = _RAND_439[7:0];
  _RAND_440 = {1{`RANDOM}};
  lineBuffer_433 = _RAND_440[7:0];
  _RAND_441 = {1{`RANDOM}};
  lineBuffer_434 = _RAND_441[7:0];
  _RAND_442 = {1{`RANDOM}};
  lineBuffer_435 = _RAND_442[7:0];
  _RAND_443 = {1{`RANDOM}};
  lineBuffer_436 = _RAND_443[7:0];
  _RAND_444 = {1{`RANDOM}};
  lineBuffer_437 = _RAND_444[7:0];
  _RAND_445 = {1{`RANDOM}};
  lineBuffer_438 = _RAND_445[7:0];
  _RAND_446 = {1{`RANDOM}};
  lineBuffer_439 = _RAND_446[7:0];
  _RAND_447 = {1{`RANDOM}};
  lineBuffer_440 = _RAND_447[7:0];
  _RAND_448 = {1{`RANDOM}};
  lineBuffer_441 = _RAND_448[7:0];
  _RAND_449 = {1{`RANDOM}};
  lineBuffer_442 = _RAND_449[7:0];
  _RAND_450 = {1{`RANDOM}};
  lineBuffer_443 = _RAND_450[7:0];
  _RAND_451 = {1{`RANDOM}};
  lineBuffer_444 = _RAND_451[7:0];
  _RAND_452 = {1{`RANDOM}};
  lineBuffer_445 = _RAND_452[7:0];
  _RAND_453 = {1{`RANDOM}};
  lineBuffer_446 = _RAND_453[7:0];
  _RAND_454 = {1{`RANDOM}};
  lineBuffer_447 = _RAND_454[7:0];
  _RAND_455 = {1{`RANDOM}};
  lineBuffer_448 = _RAND_455[7:0];
  _RAND_456 = {1{`RANDOM}};
  lineBuffer_449 = _RAND_456[7:0];
  _RAND_457 = {1{`RANDOM}};
  lineBuffer_450 = _RAND_457[7:0];
  _RAND_458 = {1{`RANDOM}};
  lineBuffer_451 = _RAND_458[7:0];
  _RAND_459 = {1{`RANDOM}};
  lineBuffer_452 = _RAND_459[7:0];
  _RAND_460 = {1{`RANDOM}};
  lineBuffer_453 = _RAND_460[7:0];
  _RAND_461 = {1{`RANDOM}};
  lineBuffer_454 = _RAND_461[7:0];
  _RAND_462 = {1{`RANDOM}};
  lineBuffer_455 = _RAND_462[7:0];
  _RAND_463 = {1{`RANDOM}};
  lineBuffer_456 = _RAND_463[7:0];
  _RAND_464 = {1{`RANDOM}};
  lineBuffer_457 = _RAND_464[7:0];
  _RAND_465 = {1{`RANDOM}};
  lineBuffer_458 = _RAND_465[7:0];
  _RAND_466 = {1{`RANDOM}};
  lineBuffer_459 = _RAND_466[7:0];
  _RAND_467 = {1{`RANDOM}};
  lineBuffer_460 = _RAND_467[7:0];
  _RAND_468 = {1{`RANDOM}};
  lineBuffer_461 = _RAND_468[7:0];
  _RAND_469 = {1{`RANDOM}};
  lineBuffer_462 = _RAND_469[7:0];
  _RAND_470 = {1{`RANDOM}};
  lineBuffer_463 = _RAND_470[7:0];
  _RAND_471 = {1{`RANDOM}};
  lineBuffer_464 = _RAND_471[7:0];
  _RAND_472 = {1{`RANDOM}};
  lineBuffer_465 = _RAND_472[7:0];
  _RAND_473 = {1{`RANDOM}};
  lineBuffer_466 = _RAND_473[7:0];
  _RAND_474 = {1{`RANDOM}};
  lineBuffer_467 = _RAND_474[7:0];
  _RAND_475 = {1{`RANDOM}};
  lineBuffer_468 = _RAND_475[7:0];
  _RAND_476 = {1{`RANDOM}};
  lineBuffer_469 = _RAND_476[7:0];
  _RAND_477 = {1{`RANDOM}};
  lineBuffer_470 = _RAND_477[7:0];
  _RAND_478 = {1{`RANDOM}};
  lineBuffer_471 = _RAND_478[7:0];
  _RAND_479 = {1{`RANDOM}};
  lineBuffer_472 = _RAND_479[7:0];
  _RAND_480 = {1{`RANDOM}};
  lineBuffer_473 = _RAND_480[7:0];
  _RAND_481 = {1{`RANDOM}};
  lineBuffer_474 = _RAND_481[7:0];
  _RAND_482 = {1{`RANDOM}};
  lineBuffer_475 = _RAND_482[7:0];
  _RAND_483 = {1{`RANDOM}};
  lineBuffer_476 = _RAND_483[7:0];
  _RAND_484 = {1{`RANDOM}};
  lineBuffer_477 = _RAND_484[7:0];
  _RAND_485 = {1{`RANDOM}};
  lineBuffer_478 = _RAND_485[7:0];
  _RAND_486 = {1{`RANDOM}};
  lineBuffer_479 = _RAND_486[7:0];
  _RAND_487 = {1{`RANDOM}};
  lineBuffer_480 = _RAND_487[7:0];
  _RAND_488 = {1{`RANDOM}};
  lineBuffer_481 = _RAND_488[7:0];
  _RAND_489 = {1{`RANDOM}};
  lineBuffer_482 = _RAND_489[7:0];
  _RAND_490 = {1{`RANDOM}};
  lineBuffer_483 = _RAND_490[7:0];
  _RAND_491 = {1{`RANDOM}};
  lineBuffer_484 = _RAND_491[7:0];
  _RAND_492 = {1{`RANDOM}};
  lineBuffer_485 = _RAND_492[7:0];
  _RAND_493 = {1{`RANDOM}};
  lineBuffer_486 = _RAND_493[7:0];
  _RAND_494 = {1{`RANDOM}};
  lineBuffer_487 = _RAND_494[7:0];
  _RAND_495 = {1{`RANDOM}};
  lineBuffer_488 = _RAND_495[7:0];
  _RAND_496 = {1{`RANDOM}};
  lineBuffer_489 = _RAND_496[7:0];
  _RAND_497 = {1{`RANDOM}};
  lineBuffer_490 = _RAND_497[7:0];
  _RAND_498 = {1{`RANDOM}};
  lineBuffer_491 = _RAND_498[7:0];
  _RAND_499 = {1{`RANDOM}};
  lineBuffer_492 = _RAND_499[7:0];
  _RAND_500 = {1{`RANDOM}};
  lineBuffer_493 = _RAND_500[7:0];
  _RAND_501 = {1{`RANDOM}};
  lineBuffer_494 = _RAND_501[7:0];
  _RAND_502 = {1{`RANDOM}};
  lineBuffer_495 = _RAND_502[7:0];
  _RAND_503 = {1{`RANDOM}};
  lineBuffer_496 = _RAND_503[7:0];
  _RAND_504 = {1{`RANDOM}};
  lineBuffer_497 = _RAND_504[7:0];
  _RAND_505 = {1{`RANDOM}};
  lineBuffer_498 = _RAND_505[7:0];
  _RAND_506 = {1{`RANDOM}};
  lineBuffer_499 = _RAND_506[7:0];
  _RAND_507 = {1{`RANDOM}};
  lineBuffer_500 = _RAND_507[7:0];
  _RAND_508 = {1{`RANDOM}};
  lineBuffer_501 = _RAND_508[7:0];
  _RAND_509 = {1{`RANDOM}};
  lineBuffer_502 = _RAND_509[7:0];
  _RAND_510 = {1{`RANDOM}};
  lineBuffer_503 = _RAND_510[7:0];
  _RAND_511 = {1{`RANDOM}};
  lineBuffer_504 = _RAND_511[7:0];
  _RAND_512 = {1{`RANDOM}};
  lineBuffer_505 = _RAND_512[7:0];
  _RAND_513 = {1{`RANDOM}};
  lineBuffer_506 = _RAND_513[7:0];
  _RAND_514 = {1{`RANDOM}};
  lineBuffer_507 = _RAND_514[7:0];
  _RAND_515 = {1{`RANDOM}};
  lineBuffer_508 = _RAND_515[7:0];
  _RAND_516 = {1{`RANDOM}};
  lineBuffer_509 = _RAND_516[7:0];
  _RAND_517 = {1{`RANDOM}};
  lineBuffer_510 = _RAND_517[7:0];
  _RAND_518 = {1{`RANDOM}};
  lineBuffer_511 = _RAND_518[7:0];
  _RAND_519 = {1{`RANDOM}};
  lineBuffer_512 = _RAND_519[7:0];
  _RAND_520 = {1{`RANDOM}};
  lineBuffer_513 = _RAND_520[7:0];
  _RAND_521 = {1{`RANDOM}};
  lineBuffer_514 = _RAND_521[7:0];
  _RAND_522 = {1{`RANDOM}};
  lineBuffer_515 = _RAND_522[7:0];
  _RAND_523 = {1{`RANDOM}};
  lineBuffer_516 = _RAND_523[7:0];
  _RAND_524 = {1{`RANDOM}};
  lineBuffer_517 = _RAND_524[7:0];
  _RAND_525 = {1{`RANDOM}};
  lineBuffer_518 = _RAND_525[7:0];
  _RAND_526 = {1{`RANDOM}};
  lineBuffer_519 = _RAND_526[7:0];
  _RAND_527 = {1{`RANDOM}};
  lineBuffer_520 = _RAND_527[7:0];
  _RAND_528 = {1{`RANDOM}};
  lineBuffer_521 = _RAND_528[7:0];
  _RAND_529 = {1{`RANDOM}};
  lineBuffer_522 = _RAND_529[7:0];
  _RAND_530 = {1{`RANDOM}};
  lineBuffer_523 = _RAND_530[7:0];
  _RAND_531 = {1{`RANDOM}};
  lineBuffer_524 = _RAND_531[7:0];
  _RAND_532 = {1{`RANDOM}};
  lineBuffer_525 = _RAND_532[7:0];
  _RAND_533 = {1{`RANDOM}};
  lineBuffer_526 = _RAND_533[7:0];
  _RAND_534 = {1{`RANDOM}};
  lineBuffer_527 = _RAND_534[7:0];
  _RAND_535 = {1{`RANDOM}};
  lineBuffer_528 = _RAND_535[7:0];
  _RAND_536 = {1{`RANDOM}};
  lineBuffer_529 = _RAND_536[7:0];
  _RAND_537 = {1{`RANDOM}};
  lineBuffer_530 = _RAND_537[7:0];
  _RAND_538 = {1{`RANDOM}};
  lineBuffer_531 = _RAND_538[7:0];
  _RAND_539 = {1{`RANDOM}};
  lineBuffer_532 = _RAND_539[7:0];
  _RAND_540 = {1{`RANDOM}};
  lineBuffer_533 = _RAND_540[7:0];
  _RAND_541 = {1{`RANDOM}};
  lineBuffer_534 = _RAND_541[7:0];
  _RAND_542 = {1{`RANDOM}};
  lineBuffer_535 = _RAND_542[7:0];
  _RAND_543 = {1{`RANDOM}};
  lineBuffer_536 = _RAND_543[7:0];
  _RAND_544 = {1{`RANDOM}};
  lineBuffer_537 = _RAND_544[7:0];
  _RAND_545 = {1{`RANDOM}};
  lineBuffer_538 = _RAND_545[7:0];
  _RAND_546 = {1{`RANDOM}};
  lineBuffer_539 = _RAND_546[7:0];
  _RAND_547 = {1{`RANDOM}};
  lineBuffer_540 = _RAND_547[7:0];
  _RAND_548 = {1{`RANDOM}};
  lineBuffer_541 = _RAND_548[7:0];
  _RAND_549 = {1{`RANDOM}};
  lineBuffer_542 = _RAND_549[7:0];
  _RAND_550 = {1{`RANDOM}};
  lineBuffer_543 = _RAND_550[7:0];
  _RAND_551 = {1{`RANDOM}};
  lineBuffer_544 = _RAND_551[7:0];
  _RAND_552 = {1{`RANDOM}};
  lineBuffer_545 = _RAND_552[7:0];
  _RAND_553 = {1{`RANDOM}};
  lineBuffer_546 = _RAND_553[7:0];
  _RAND_554 = {1{`RANDOM}};
  lineBuffer_547 = _RAND_554[7:0];
  _RAND_555 = {1{`RANDOM}};
  lineBuffer_548 = _RAND_555[7:0];
  _RAND_556 = {1{`RANDOM}};
  lineBuffer_549 = _RAND_556[7:0];
  _RAND_557 = {1{`RANDOM}};
  lineBuffer_550 = _RAND_557[7:0];
  _RAND_558 = {1{`RANDOM}};
  lineBuffer_551 = _RAND_558[7:0];
  _RAND_559 = {1{`RANDOM}};
  lineBuffer_552 = _RAND_559[7:0];
  _RAND_560 = {1{`RANDOM}};
  lineBuffer_553 = _RAND_560[7:0];
  _RAND_561 = {1{`RANDOM}};
  lineBuffer_554 = _RAND_561[7:0];
  _RAND_562 = {1{`RANDOM}};
  lineBuffer_555 = _RAND_562[7:0];
  _RAND_563 = {1{`RANDOM}};
  lineBuffer_556 = _RAND_563[7:0];
  _RAND_564 = {1{`RANDOM}};
  lineBuffer_557 = _RAND_564[7:0];
  _RAND_565 = {1{`RANDOM}};
  lineBuffer_558 = _RAND_565[7:0];
  _RAND_566 = {1{`RANDOM}};
  lineBuffer_559 = _RAND_566[7:0];
  _RAND_567 = {1{`RANDOM}};
  lineBuffer_560 = _RAND_567[7:0];
  _RAND_568 = {1{`RANDOM}};
  lineBuffer_561 = _RAND_568[7:0];
  _RAND_569 = {1{`RANDOM}};
  lineBuffer_562 = _RAND_569[7:0];
  _RAND_570 = {1{`RANDOM}};
  lineBuffer_563 = _RAND_570[7:0];
  _RAND_571 = {1{`RANDOM}};
  lineBuffer_564 = _RAND_571[7:0];
  _RAND_572 = {1{`RANDOM}};
  lineBuffer_565 = _RAND_572[7:0];
  _RAND_573 = {1{`RANDOM}};
  lineBuffer_566 = _RAND_573[7:0];
  _RAND_574 = {1{`RANDOM}};
  lineBuffer_567 = _RAND_574[7:0];
  _RAND_575 = {1{`RANDOM}};
  lineBuffer_568 = _RAND_575[7:0];
  _RAND_576 = {1{`RANDOM}};
  lineBuffer_569 = _RAND_576[7:0];
  _RAND_577 = {1{`RANDOM}};
  lineBuffer_570 = _RAND_577[7:0];
  _RAND_578 = {1{`RANDOM}};
  lineBuffer_571 = _RAND_578[7:0];
  _RAND_579 = {1{`RANDOM}};
  lineBuffer_572 = _RAND_579[7:0];
  _RAND_580 = {1{`RANDOM}};
  lineBuffer_573 = _RAND_580[7:0];
  _RAND_581 = {1{`RANDOM}};
  lineBuffer_574 = _RAND_581[7:0];
  _RAND_582 = {1{`RANDOM}};
  lineBuffer_575 = _RAND_582[7:0];
  _RAND_583 = {1{`RANDOM}};
  lineBuffer_576 = _RAND_583[7:0];
  _RAND_584 = {1{`RANDOM}};
  lineBuffer_577 = _RAND_584[7:0];
  _RAND_585 = {1{`RANDOM}};
  lineBuffer_578 = _RAND_585[7:0];
  _RAND_586 = {1{`RANDOM}};
  lineBuffer_579 = _RAND_586[7:0];
  _RAND_587 = {1{`RANDOM}};
  lineBuffer_580 = _RAND_587[7:0];
  _RAND_588 = {1{`RANDOM}};
  lineBuffer_581 = _RAND_588[7:0];
  _RAND_589 = {1{`RANDOM}};
  lineBuffer_582 = _RAND_589[7:0];
  _RAND_590 = {1{`RANDOM}};
  lineBuffer_583 = _RAND_590[7:0];
  _RAND_591 = {1{`RANDOM}};
  lineBuffer_584 = _RAND_591[7:0];
  _RAND_592 = {1{`RANDOM}};
  lineBuffer_585 = _RAND_592[7:0];
  _RAND_593 = {1{`RANDOM}};
  lineBuffer_586 = _RAND_593[7:0];
  _RAND_594 = {1{`RANDOM}};
  lineBuffer_587 = _RAND_594[7:0];
  _RAND_595 = {1{`RANDOM}};
  lineBuffer_588 = _RAND_595[7:0];
  _RAND_596 = {1{`RANDOM}};
  lineBuffer_589 = _RAND_596[7:0];
  _RAND_597 = {1{`RANDOM}};
  lineBuffer_590 = _RAND_597[7:0];
  _RAND_598 = {1{`RANDOM}};
  lineBuffer_591 = _RAND_598[7:0];
  _RAND_599 = {1{`RANDOM}};
  lineBuffer_592 = _RAND_599[7:0];
  _RAND_600 = {1{`RANDOM}};
  lineBuffer_593 = _RAND_600[7:0];
  _RAND_601 = {1{`RANDOM}};
  lineBuffer_594 = _RAND_601[7:0];
  _RAND_602 = {1{`RANDOM}};
  lineBuffer_595 = _RAND_602[7:0];
  _RAND_603 = {1{`RANDOM}};
  lineBuffer_596 = _RAND_603[7:0];
  _RAND_604 = {1{`RANDOM}};
  lineBuffer_597 = _RAND_604[7:0];
  _RAND_605 = {1{`RANDOM}};
  lineBuffer_598 = _RAND_605[7:0];
  _RAND_606 = {1{`RANDOM}};
  lineBuffer_599 = _RAND_606[7:0];
  _RAND_607 = {1{`RANDOM}};
  lineBuffer_600 = _RAND_607[7:0];
  _RAND_608 = {1{`RANDOM}};
  lineBuffer_601 = _RAND_608[7:0];
  _RAND_609 = {1{`RANDOM}};
  lineBuffer_602 = _RAND_609[7:0];
  _RAND_610 = {1{`RANDOM}};
  lineBuffer_603 = _RAND_610[7:0];
  _RAND_611 = {1{`RANDOM}};
  lineBuffer_604 = _RAND_611[7:0];
  _RAND_612 = {1{`RANDOM}};
  lineBuffer_605 = _RAND_612[7:0];
  _RAND_613 = {1{`RANDOM}};
  lineBuffer_606 = _RAND_613[7:0];
  _RAND_614 = {1{`RANDOM}};
  lineBuffer_607 = _RAND_614[7:0];
  _RAND_615 = {1{`RANDOM}};
  lineBuffer_608 = _RAND_615[7:0];
  _RAND_616 = {1{`RANDOM}};
  lineBuffer_609 = _RAND_616[7:0];
  _RAND_617 = {1{`RANDOM}};
  lineBuffer_610 = _RAND_617[7:0];
  _RAND_618 = {1{`RANDOM}};
  lineBuffer_611 = _RAND_618[7:0];
  _RAND_619 = {1{`RANDOM}};
  lineBuffer_612 = _RAND_619[7:0];
  _RAND_620 = {1{`RANDOM}};
  lineBuffer_613 = _RAND_620[7:0];
  _RAND_621 = {1{`RANDOM}};
  lineBuffer_614 = _RAND_621[7:0];
  _RAND_622 = {1{`RANDOM}};
  lineBuffer_615 = _RAND_622[7:0];
  _RAND_623 = {1{`RANDOM}};
  lineBuffer_616 = _RAND_623[7:0];
  _RAND_624 = {1{`RANDOM}};
  lineBuffer_617 = _RAND_624[7:0];
  _RAND_625 = {1{`RANDOM}};
  lineBuffer_618 = _RAND_625[7:0];
  _RAND_626 = {1{`RANDOM}};
  lineBuffer_619 = _RAND_626[7:0];
  _RAND_627 = {1{`RANDOM}};
  lineBuffer_620 = _RAND_627[7:0];
  _RAND_628 = {1{`RANDOM}};
  lineBuffer_621 = _RAND_628[7:0];
  _RAND_629 = {1{`RANDOM}};
  lineBuffer_622 = _RAND_629[7:0];
  _RAND_630 = {1{`RANDOM}};
  lineBuffer_623 = _RAND_630[7:0];
  _RAND_631 = {1{`RANDOM}};
  lineBuffer_624 = _RAND_631[7:0];
  _RAND_632 = {1{`RANDOM}};
  lineBuffer_625 = _RAND_632[7:0];
  _RAND_633 = {1{`RANDOM}};
  lineBuffer_626 = _RAND_633[7:0];
  _RAND_634 = {1{`RANDOM}};
  lineBuffer_627 = _RAND_634[7:0];
  _RAND_635 = {1{`RANDOM}};
  lineBuffer_628 = _RAND_635[7:0];
  _RAND_636 = {1{`RANDOM}};
  lineBuffer_629 = _RAND_636[7:0];
  _RAND_637 = {1{`RANDOM}};
  lineBuffer_630 = _RAND_637[7:0];
  _RAND_638 = {1{`RANDOM}};
  lineBuffer_631 = _RAND_638[7:0];
  _RAND_639 = {1{`RANDOM}};
  lineBuffer_632 = _RAND_639[7:0];
  _RAND_640 = {1{`RANDOM}};
  lineBuffer_633 = _RAND_640[7:0];
  _RAND_641 = {1{`RANDOM}};
  lineBuffer_634 = _RAND_641[7:0];
  _RAND_642 = {1{`RANDOM}};
  lineBuffer_635 = _RAND_642[7:0];
  _RAND_643 = {1{`RANDOM}};
  lineBuffer_636 = _RAND_643[7:0];
  _RAND_644 = {1{`RANDOM}};
  lineBuffer_637 = _RAND_644[7:0];
  _RAND_645 = {1{`RANDOM}};
  lineBuffer_638 = _RAND_645[7:0];
  _RAND_646 = {1{`RANDOM}};
  lineBuffer_639 = _RAND_646[7:0];
  _RAND_647 = {1{`RANDOM}};
  lineBuffer_640 = _RAND_647[7:0];
  _RAND_648 = {1{`RANDOM}};
  lineBuffer_641 = _RAND_648[7:0];
  _RAND_649 = {1{`RANDOM}};
  lineBuffer_642 = _RAND_649[7:0];
  _RAND_650 = {1{`RANDOM}};
  lineBuffer_643 = _RAND_650[7:0];
  _RAND_651 = {1{`RANDOM}};
  lineBuffer_644 = _RAND_651[7:0];
  _RAND_652 = {1{`RANDOM}};
  lineBuffer_645 = _RAND_652[7:0];
  _RAND_653 = {1{`RANDOM}};
  lineBuffer_646 = _RAND_653[7:0];
  _RAND_654 = {1{`RANDOM}};
  lineBuffer_647 = _RAND_654[7:0];
  _RAND_655 = {1{`RANDOM}};
  lineBuffer_648 = _RAND_655[7:0];
  _RAND_656 = {1{`RANDOM}};
  lineBuffer_649 = _RAND_656[7:0];
  _RAND_657 = {1{`RANDOM}};
  lineBuffer_650 = _RAND_657[7:0];
  _RAND_658 = {1{`RANDOM}};
  lineBuffer_651 = _RAND_658[7:0];
  _RAND_659 = {1{`RANDOM}};
  lineBuffer_652 = _RAND_659[7:0];
  _RAND_660 = {1{`RANDOM}};
  lineBuffer_653 = _RAND_660[7:0];
  _RAND_661 = {1{`RANDOM}};
  lineBuffer_654 = _RAND_661[7:0];
  _RAND_662 = {1{`RANDOM}};
  lineBuffer_655 = _RAND_662[7:0];
  _RAND_663 = {1{`RANDOM}};
  lineBuffer_656 = _RAND_663[7:0];
  _RAND_664 = {1{`RANDOM}};
  lineBuffer_657 = _RAND_664[7:0];
  _RAND_665 = {1{`RANDOM}};
  lineBuffer_658 = _RAND_665[7:0];
  _RAND_666 = {1{`RANDOM}};
  lineBuffer_659 = _RAND_666[7:0];
  _RAND_667 = {1{`RANDOM}};
  lineBuffer_660 = _RAND_667[7:0];
  _RAND_668 = {1{`RANDOM}};
  lineBuffer_661 = _RAND_668[7:0];
  _RAND_669 = {1{`RANDOM}};
  lineBuffer_662 = _RAND_669[7:0];
  _RAND_670 = {1{`RANDOM}};
  lineBuffer_663 = _RAND_670[7:0];
  _RAND_671 = {1{`RANDOM}};
  lineBuffer_664 = _RAND_671[7:0];
  _RAND_672 = {1{`RANDOM}};
  lineBuffer_665 = _RAND_672[7:0];
  _RAND_673 = {1{`RANDOM}};
  lineBuffer_666 = _RAND_673[7:0];
  _RAND_674 = {1{`RANDOM}};
  lineBuffer_667 = _RAND_674[7:0];
  _RAND_675 = {1{`RANDOM}};
  lineBuffer_668 = _RAND_675[7:0];
  _RAND_676 = {1{`RANDOM}};
  lineBuffer_669 = _RAND_676[7:0];
  _RAND_677 = {1{`RANDOM}};
  lineBuffer_670 = _RAND_677[7:0];
  _RAND_678 = {1{`RANDOM}};
  lineBuffer_671 = _RAND_678[7:0];
  _RAND_679 = {1{`RANDOM}};
  lineBuffer_672 = _RAND_679[7:0];
  _RAND_680 = {1{`RANDOM}};
  lineBuffer_673 = _RAND_680[7:0];
  _RAND_681 = {1{`RANDOM}};
  lineBuffer_674 = _RAND_681[7:0];
  _RAND_682 = {1{`RANDOM}};
  lineBuffer_675 = _RAND_682[7:0];
  _RAND_683 = {1{`RANDOM}};
  lineBuffer_676 = _RAND_683[7:0];
  _RAND_684 = {1{`RANDOM}};
  lineBuffer_677 = _RAND_684[7:0];
  _RAND_685 = {1{`RANDOM}};
  lineBuffer_678 = _RAND_685[7:0];
  _RAND_686 = {1{`RANDOM}};
  lineBuffer_679 = _RAND_686[7:0];
  _RAND_687 = {1{`RANDOM}};
  lineBuffer_680 = _RAND_687[7:0];
  _RAND_688 = {1{`RANDOM}};
  lineBuffer_681 = _RAND_688[7:0];
  _RAND_689 = {1{`RANDOM}};
  lineBuffer_682 = _RAND_689[7:0];
  _RAND_690 = {1{`RANDOM}};
  lineBuffer_683 = _RAND_690[7:0];
  _RAND_691 = {1{`RANDOM}};
  lineBuffer_684 = _RAND_691[7:0];
  _RAND_692 = {1{`RANDOM}};
  lineBuffer_685 = _RAND_692[7:0];
  _RAND_693 = {1{`RANDOM}};
  lineBuffer_686 = _RAND_693[7:0];
  _RAND_694 = {1{`RANDOM}};
  lineBuffer_687 = _RAND_694[7:0];
  _RAND_695 = {1{`RANDOM}};
  lineBuffer_688 = _RAND_695[7:0];
  _RAND_696 = {1{`RANDOM}};
  lineBuffer_689 = _RAND_696[7:0];
  _RAND_697 = {1{`RANDOM}};
  lineBuffer_690 = _RAND_697[7:0];
  _RAND_698 = {1{`RANDOM}};
  lineBuffer_691 = _RAND_698[7:0];
  _RAND_699 = {1{`RANDOM}};
  lineBuffer_692 = _RAND_699[7:0];
  _RAND_700 = {1{`RANDOM}};
  lineBuffer_693 = _RAND_700[7:0];
  _RAND_701 = {1{`RANDOM}};
  lineBuffer_694 = _RAND_701[7:0];
  _RAND_702 = {1{`RANDOM}};
  lineBuffer_695 = _RAND_702[7:0];
  _RAND_703 = {1{`RANDOM}};
  lineBuffer_696 = _RAND_703[7:0];
  _RAND_704 = {1{`RANDOM}};
  lineBuffer_697 = _RAND_704[7:0];
  _RAND_705 = {1{`RANDOM}};
  lineBuffer_698 = _RAND_705[7:0];
  _RAND_706 = {1{`RANDOM}};
  lineBuffer_699 = _RAND_706[7:0];
  _RAND_707 = {1{`RANDOM}};
  lineBuffer_700 = _RAND_707[7:0];
  _RAND_708 = {1{`RANDOM}};
  lineBuffer_701 = _RAND_708[7:0];
  _RAND_709 = {1{`RANDOM}};
  lineBuffer_702 = _RAND_709[7:0];
  _RAND_710 = {1{`RANDOM}};
  lineBuffer_703 = _RAND_710[7:0];
  _RAND_711 = {1{`RANDOM}};
  lineBuffer_704 = _RAND_711[7:0];
  _RAND_712 = {1{`RANDOM}};
  lineBuffer_705 = _RAND_712[7:0];
  _RAND_713 = {1{`RANDOM}};
  lineBuffer_706 = _RAND_713[7:0];
  _RAND_714 = {1{`RANDOM}};
  lineBuffer_707 = _RAND_714[7:0];
  _RAND_715 = {1{`RANDOM}};
  lineBuffer_708 = _RAND_715[7:0];
  _RAND_716 = {1{`RANDOM}};
  lineBuffer_709 = _RAND_716[7:0];
  _RAND_717 = {1{`RANDOM}};
  lineBuffer_710 = _RAND_717[7:0];
  _RAND_718 = {1{`RANDOM}};
  lineBuffer_711 = _RAND_718[7:0];
  _RAND_719 = {1{`RANDOM}};
  lineBuffer_712 = _RAND_719[7:0];
  _RAND_720 = {1{`RANDOM}};
  lineBuffer_713 = _RAND_720[7:0];
  _RAND_721 = {1{`RANDOM}};
  lineBuffer_714 = _RAND_721[7:0];
  _RAND_722 = {1{`RANDOM}};
  lineBuffer_715 = _RAND_722[7:0];
  _RAND_723 = {1{`RANDOM}};
  lineBuffer_716 = _RAND_723[7:0];
  _RAND_724 = {1{`RANDOM}};
  lineBuffer_717 = _RAND_724[7:0];
  _RAND_725 = {1{`RANDOM}};
  lineBuffer_718 = _RAND_725[7:0];
  _RAND_726 = {1{`RANDOM}};
  lineBuffer_719 = _RAND_726[7:0];
  _RAND_727 = {1{`RANDOM}};
  lineBuffer_720 = _RAND_727[7:0];
  _RAND_728 = {1{`RANDOM}};
  lineBuffer_721 = _RAND_728[7:0];
  _RAND_729 = {1{`RANDOM}};
  lineBuffer_722 = _RAND_729[7:0];
  _RAND_730 = {1{`RANDOM}};
  lineBuffer_723 = _RAND_730[7:0];
  _RAND_731 = {1{`RANDOM}};
  lineBuffer_724 = _RAND_731[7:0];
  _RAND_732 = {1{`RANDOM}};
  lineBuffer_725 = _RAND_732[7:0];
  _RAND_733 = {1{`RANDOM}};
  lineBuffer_726 = _RAND_733[7:0];
  _RAND_734 = {1{`RANDOM}};
  lineBuffer_727 = _RAND_734[7:0];
  _RAND_735 = {1{`RANDOM}};
  lineBuffer_728 = _RAND_735[7:0];
  _RAND_736 = {1{`RANDOM}};
  lineBuffer_729 = _RAND_736[7:0];
  _RAND_737 = {1{`RANDOM}};
  lineBuffer_730 = _RAND_737[7:0];
  _RAND_738 = {1{`RANDOM}};
  lineBuffer_731 = _RAND_738[7:0];
  _RAND_739 = {1{`RANDOM}};
  lineBuffer_732 = _RAND_739[7:0];
  _RAND_740 = {1{`RANDOM}};
  lineBuffer_733 = _RAND_740[7:0];
  _RAND_741 = {1{`RANDOM}};
  lineBuffer_734 = _RAND_741[7:0];
  _RAND_742 = {1{`RANDOM}};
  lineBuffer_735 = _RAND_742[7:0];
  _RAND_743 = {1{`RANDOM}};
  lineBuffer_736 = _RAND_743[7:0];
  _RAND_744 = {1{`RANDOM}};
  lineBuffer_737 = _RAND_744[7:0];
  _RAND_745 = {1{`RANDOM}};
  lineBuffer_738 = _RAND_745[7:0];
  _RAND_746 = {1{`RANDOM}};
  lineBuffer_739 = _RAND_746[7:0];
  _RAND_747 = {1{`RANDOM}};
  lineBuffer_740 = _RAND_747[7:0];
  _RAND_748 = {1{`RANDOM}};
  lineBuffer_741 = _RAND_748[7:0];
  _RAND_749 = {1{`RANDOM}};
  lineBuffer_742 = _RAND_749[7:0];
  _RAND_750 = {1{`RANDOM}};
  lineBuffer_743 = _RAND_750[7:0];
  _RAND_751 = {1{`RANDOM}};
  lineBuffer_744 = _RAND_751[7:0];
  _RAND_752 = {1{`RANDOM}};
  lineBuffer_745 = _RAND_752[7:0];
  _RAND_753 = {1{`RANDOM}};
  lineBuffer_746 = _RAND_753[7:0];
  _RAND_754 = {1{`RANDOM}};
  lineBuffer_747 = _RAND_754[7:0];
  _RAND_755 = {1{`RANDOM}};
  lineBuffer_748 = _RAND_755[7:0];
  _RAND_756 = {1{`RANDOM}};
  lineBuffer_749 = _RAND_756[7:0];
  _RAND_757 = {1{`RANDOM}};
  lineBuffer_750 = _RAND_757[7:0];
  _RAND_758 = {1{`RANDOM}};
  lineBuffer_751 = _RAND_758[7:0];
  _RAND_759 = {1{`RANDOM}};
  lineBuffer_752 = _RAND_759[7:0];
  _RAND_760 = {1{`RANDOM}};
  lineBuffer_753 = _RAND_760[7:0];
  _RAND_761 = {1{`RANDOM}};
  lineBuffer_754 = _RAND_761[7:0];
  _RAND_762 = {1{`RANDOM}};
  lineBuffer_755 = _RAND_762[7:0];
  _RAND_763 = {1{`RANDOM}};
  lineBuffer_756 = _RAND_763[7:0];
  _RAND_764 = {1{`RANDOM}};
  lineBuffer_757 = _RAND_764[7:0];
  _RAND_765 = {1{`RANDOM}};
  lineBuffer_758 = _RAND_765[7:0];
  _RAND_766 = {1{`RANDOM}};
  lineBuffer_759 = _RAND_766[7:0];
  _RAND_767 = {1{`RANDOM}};
  lineBuffer_760 = _RAND_767[7:0];
  _RAND_768 = {1{`RANDOM}};
  lineBuffer_761 = _RAND_768[7:0];
  _RAND_769 = {1{`RANDOM}};
  lineBuffer_762 = _RAND_769[7:0];
  _RAND_770 = {1{`RANDOM}};
  lineBuffer_763 = _RAND_770[7:0];
  _RAND_771 = {1{`RANDOM}};
  lineBuffer_764 = _RAND_771[7:0];
  _RAND_772 = {1{`RANDOM}};
  lineBuffer_765 = _RAND_772[7:0];
  _RAND_773 = {1{`RANDOM}};
  lineBuffer_766 = _RAND_773[7:0];
  _RAND_774 = {1{`RANDOM}};
  lineBuffer_767 = _RAND_774[7:0];
  _RAND_775 = {1{`RANDOM}};
  windowBuffer_0 = _RAND_775[7:0];
  _RAND_776 = {1{`RANDOM}};
  windowBuffer_1 = _RAND_776[7:0];
  _RAND_777 = {1{`RANDOM}};
  windowBuffer_2 = _RAND_777[7:0];
  _RAND_778 = {1{`RANDOM}};
  windowBuffer_3 = _RAND_778[7:0];
  _RAND_779 = {1{`RANDOM}};
  windowBuffer_4 = _RAND_779[7:0];
  _RAND_780 = {1{`RANDOM}};
  windowBuffer_5 = _RAND_780[7:0];
  _RAND_781 = {1{`RANDOM}};
  windowBuffer_6 = _RAND_781[7:0];
  _RAND_782 = {1{`RANDOM}};
  windowBuffer_7 = _RAND_782[7:0];
  _RAND_783 = {1{`RANDOM}};
  windowBuffer_8 = _RAND_783[7:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      stateReg <= 2'h0;
    end else if (_T) begin
      if (io_enq_valid) begin
        stateReg <= 2'h1;
      end else if (_T) begin
        if (io_enq_valid) begin
          stateReg <= 2'h1;
        end
      end else if (_T_1) begin
        if (_T_3) begin
          stateReg <= 2'h0;
        end else if (_T_4) begin
          stateReg <= 2'h1;
        end else if (_T_6) begin
          stateReg <= 2'h2;
        end
      end else if (_T_7) begin
        if (io_deq_ready) begin
          stateReg <= 2'h1;
        end
      end else if (_T_8) begin
        stateReg <= 2'h0;
      end
    end else if (_T_1) begin
      if (_T_3) begin
        stateReg <= 2'h0;
      end else if (_T_4) begin
        stateReg <= 2'h1;
      end else if (_T_6) begin
        stateReg <= 2'h2;
      end else if (_T) begin
        if (io_enq_valid) begin
          stateReg <= 2'h1;
        end
      end else if (_T_1) begin
        if (_T_3) begin
          stateReg <= 2'h0;
        end else if (_T_4) begin
          stateReg <= 2'h1;
        end else if (_T_6) begin
          stateReg <= 2'h2;
        end
      end else if (_T_7) begin
        if (io_deq_ready) begin
          stateReg <= 2'h1;
        end
      end else if (_T_8) begin
        stateReg <= 2'h0;
      end
    end else if (_T_7) begin
      if (io_deq_ready) begin
        stateReg <= 2'h1;
      end else if (_T) begin
        if (io_enq_valid) begin
          stateReg <= 2'h1;
        end
      end else if (_T_1) begin
        if (_T_3) begin
          stateReg <= 2'h0;
        end else if (_T_4) begin
          stateReg <= 2'h1;
        end else if (_T_6) begin
          stateReg <= 2'h2;
        end
      end else if (_T_7) begin
        if (io_deq_ready) begin
          stateReg <= 2'h1;
        end
      end else if (_T_8) begin
        stateReg <= 2'h0;
      end
    end else if (_T_8) begin
      stateReg <= 2'h0;
    end else if (_T) begin
      if (io_enq_valid) begin
        stateReg <= 2'h1;
      end
    end else if (_T_1) begin
      if (_T_3) begin
        stateReg <= 2'h0;
      end else if (_T_4) begin
        stateReg <= 2'h1;
      end else if (_T_6) begin
        stateReg <= 2'h2;
      end
    end else if (_T_7) begin
      if (io_deq_ready) begin
        stateReg <= 2'h1;
      end
    end else if (_T_8) begin
      stateReg <= 2'h0;
    end
    if (_T) begin
      if (io_enq_valid) begin
        dataReg <= io_enq_bits;
      end else if (_T) begin
        if (io_enq_valid) begin
          dataReg <= io_enq_bits;
        end
      end else if (_T_1) begin
        if (!(_T_3)) begin
          if (_T_4) begin
            dataReg <= io_enq_bits;
          end
        end
      end else if (_T_7) begin
        if (io_deq_ready) begin
          dataReg <= shadowReg;
        end
      end
    end else if (_T_1) begin
      if (_T_3) begin
        if (_T) begin
          if (io_enq_valid) begin
            dataReg <= io_enq_bits;
          end
        end else if (_T_1) begin
          if (!(_T_3)) begin
            if (_T_4) begin
              dataReg <= io_enq_bits;
            end
          end
        end else if (_T_7) begin
          if (io_deq_ready) begin
            dataReg <= shadowReg;
          end
        end
      end else if (_T_4) begin
        dataReg <= io_enq_bits;
      end else if (_T) begin
        if (io_enq_valid) begin
          dataReg <= io_enq_bits;
        end
      end else if (_T_1) begin
        if (!(_T_3)) begin
          if (_T_4) begin
            dataReg <= io_enq_bits;
          end
        end
      end else if (_T_7) begin
        if (io_deq_ready) begin
          dataReg <= shadowReg;
        end
      end
    end else if (_T_7) begin
      if (io_deq_ready) begin
        dataReg <= shadowReg;
      end else if (_T) begin
        if (io_enq_valid) begin
          dataReg <= io_enq_bits;
        end
      end else if (_T_1) begin
        if (!(_T_3)) begin
          if (_T_4) begin
            dataReg <= io_enq_bits;
          end
        end
      end else if (_T_7) begin
        if (io_deq_ready) begin
          dataReg <= shadowReg;
        end
      end
    end else begin
      dataReg <= _GEN_39;
    end
    if (_T) begin
      if (!(_T)) begin
        if (_T_1) begin
          if (!(_T_3)) begin
            if (!(_T_4)) begin
              if (_T_6) begin
                shadowReg <= io_enq_bits;
              end
            end
          end
        end
      end
    end else if (_T_1) begin
      if (_T_3) begin
        if (!(_T)) begin
          if (_T_1) begin
            if (!(_T_3)) begin
              if (!(_T_4)) begin
                if (_T_6) begin
                  shadowReg <= io_enq_bits;
                end
              end
            end
          end
        end
      end else if (_T_4) begin
        if (!(_T)) begin
          if (_T_1) begin
            if (!(_T_3)) begin
              if (!(_T_4)) begin
                if (_T_6) begin
                  shadowReg <= io_enq_bits;
                end
              end
            end
          end
        end
      end else if (_T_6) begin
        shadowReg <= io_enq_bits;
      end else if (!(_T)) begin
        if (_T_1) begin
          if (!(_T_3)) begin
            if (!(_T_4)) begin
              if (_T_6) begin
                shadowReg <= io_enq_bits;
              end
            end
          end
        end
      end
    end else begin
      shadowReg <= _GEN_41;
    end
    if (_T) begin
      userReg <= io_enq_user;
    end else if (_T_1) begin
      if (_T_3) begin
        userReg <= io_enq_user;
      end else if (_T_4) begin
        userReg <= io_enq_user;
      end else if (_T) begin
        userReg <= io_enq_user;
      end else if (_T_1) begin
        if (_T_3) begin
          userReg <= io_enq_user;
        end else if (_T_4) begin
          userReg <= io_enq_user;
        end
      end else if (_T_7) begin
        if (io_deq_ready) begin
          userReg <= shadowUserReg;
        end
      end
    end else if (_T_7) begin
      if (io_deq_ready) begin
        userReg <= shadowUserReg;
      end else if (_T) begin
        userReg <= io_enq_user;
      end else if (_T_1) begin
        if (_T_3) begin
          userReg <= io_enq_user;
        end else if (_T_4) begin
          userReg <= io_enq_user;
        end
      end else if (_T_7) begin
        if (io_deq_ready) begin
          userReg <= shadowUserReg;
        end
      end
    end else if (_T) begin
      userReg <= io_enq_user;
    end else if (_T_1) begin
      if (_T_3) begin
        userReg <= io_enq_user;
      end else if (_T_4) begin
        userReg <= io_enq_user;
      end
    end else if (_T_7) begin
      if (io_deq_ready) begin
        userReg <= shadowUserReg;
      end
    end
    if (_T) begin
      if (!(_T)) begin
        if (_T_1) begin
          if (!(_T_3)) begin
            if (!(_T_4)) begin
              if (_T_6) begin
                shadowUserReg <= io_enq_user;
              end
            end
          end
        end
      end
    end else if (_T_1) begin
      if (_T_3) begin
        if (!(_T)) begin
          if (_T_1) begin
            if (!(_T_3)) begin
              if (!(_T_4)) begin
                if (_T_6) begin
                  shadowUserReg <= io_enq_user;
                end
              end
            end
          end
        end
      end else if (_T_4) begin
        if (!(_T)) begin
          if (_T_1) begin
            if (!(_T_3)) begin
              if (!(_T_4)) begin
                if (_T_6) begin
                  shadowUserReg <= io_enq_user;
                end
              end
            end
          end
        end
      end else if (_T_6) begin
        shadowUserReg <= io_enq_user;
      end else if (!(_T)) begin
        if (_T_1) begin
          if (!(_T_3)) begin
            if (!(_T_4)) begin
              if (_T_6) begin
                shadowUserReg <= io_enq_user;
              end
            end
          end
        end
      end
    end else begin
      shadowUserReg <= _GEN_42;
    end
    if (_T) begin
      if (io_enq_valid) begin
        lastReg <= io_enq_last;
      end else if (_T) begin
        if (io_enq_valid) begin
          lastReg <= io_enq_last;
        end
      end else if (_T_1) begin
        if (!(_T_3)) begin
          if (_T_4) begin
            lastReg <= io_enq_last;
          end
        end
      end else if (_T_7) begin
        if (io_deq_ready) begin
          lastReg <= shadowLastReg;
        end
      end
    end else if (_T_1) begin
      if (_T_3) begin
        if (_T) begin
          if (io_enq_valid) begin
            lastReg <= io_enq_last;
          end
        end else if (_T_1) begin
          if (!(_T_3)) begin
            if (_T_4) begin
              lastReg <= io_enq_last;
            end
          end
        end else if (_T_7) begin
          if (io_deq_ready) begin
            lastReg <= shadowLastReg;
          end
        end
      end else if (_T_4) begin
        lastReg <= io_enq_last;
      end else if (_T) begin
        if (io_enq_valid) begin
          lastReg <= io_enq_last;
        end
      end else if (_T_1) begin
        if (!(_T_3)) begin
          if (_T_4) begin
            lastReg <= io_enq_last;
          end
        end
      end else if (_T_7) begin
        if (io_deq_ready) begin
          lastReg <= shadowLastReg;
        end
      end
    end else if (_T_7) begin
      if (io_deq_ready) begin
        lastReg <= shadowLastReg;
      end else if (_T) begin
        if (io_enq_valid) begin
          lastReg <= io_enq_last;
        end
      end else if (_T_1) begin
        if (!(_T_3)) begin
          if (_T_4) begin
            lastReg <= io_enq_last;
          end
        end
      end else if (_T_7) begin
        if (io_deq_ready) begin
          lastReg <= shadowLastReg;
        end
      end
    end else begin
      lastReg <= _GEN_40;
    end
    if (_T) begin
      if (!(_T)) begin
        if (_T_1) begin
          if (!(_T_3)) begin
            if (!(_T_4)) begin
              if (_T_6) begin
                shadowLastReg <= io_enq_last;
              end
            end
          end
        end
      end
    end else if (_T_1) begin
      if (_T_3) begin
        if (!(_T)) begin
          if (_T_1) begin
            if (!(_T_3)) begin
              if (!(_T_4)) begin
                if (_T_6) begin
                  shadowLastReg <= io_enq_last;
                end
              end
            end
          end
        end
      end else if (_T_4) begin
        if (!(_T)) begin
          if (_T_1) begin
            if (!(_T_3)) begin
              if (!(_T_4)) begin
                if (_T_6) begin
                  shadowLastReg <= io_enq_last;
                end
              end
            end
          end
        end
      end else if (_T_6) begin
        shadowLastReg <= io_enq_last;
      end else if (!(_T)) begin
        if (_T_1) begin
          if (!(_T_3)) begin
            if (!(_T_4)) begin
              if (_T_6) begin
                shadowLastReg <= io_enq_last;
              end
            end
          end
        end
      end
    end else begin
      shadowLastReg <= _GEN_43;
    end
    if (sel) begin
      lineBuffer_0 <= dataReg;
    end
    if (sel) begin
      lineBuffer_1 <= lineBuffer_0;
    end
    if (sel) begin
      lineBuffer_2 <= lineBuffer_1;
    end
    if (sel) begin
      lineBuffer_3 <= lineBuffer_2;
    end
    if (sel) begin
      lineBuffer_4 <= lineBuffer_3;
    end
    if (sel) begin
      lineBuffer_5 <= lineBuffer_4;
    end
    if (sel) begin
      lineBuffer_6 <= lineBuffer_5;
    end
    if (sel) begin
      lineBuffer_7 <= lineBuffer_6;
    end
    if (sel) begin
      lineBuffer_8 <= lineBuffer_7;
    end
    if (sel) begin
      lineBuffer_9 <= lineBuffer_8;
    end
    if (sel) begin
      lineBuffer_10 <= lineBuffer_9;
    end
    if (sel) begin
      lineBuffer_11 <= lineBuffer_10;
    end
    if (sel) begin
      lineBuffer_12 <= lineBuffer_11;
    end
    if (sel) begin
      lineBuffer_13 <= lineBuffer_12;
    end
    if (sel) begin
      lineBuffer_14 <= lineBuffer_13;
    end
    if (sel) begin
      lineBuffer_15 <= lineBuffer_14;
    end
    if (sel) begin
      lineBuffer_16 <= lineBuffer_15;
    end
    if (sel) begin
      lineBuffer_17 <= lineBuffer_16;
    end
    if (sel) begin
      lineBuffer_18 <= lineBuffer_17;
    end
    if (sel) begin
      lineBuffer_19 <= lineBuffer_18;
    end
    if (sel) begin
      lineBuffer_20 <= lineBuffer_19;
    end
    if (sel) begin
      lineBuffer_21 <= lineBuffer_20;
    end
    if (sel) begin
      lineBuffer_22 <= lineBuffer_21;
    end
    if (sel) begin
      lineBuffer_23 <= lineBuffer_22;
    end
    if (sel) begin
      lineBuffer_24 <= lineBuffer_23;
    end
    if (sel) begin
      lineBuffer_25 <= lineBuffer_24;
    end
    if (sel) begin
      lineBuffer_26 <= lineBuffer_25;
    end
    if (sel) begin
      lineBuffer_27 <= lineBuffer_26;
    end
    if (sel) begin
      lineBuffer_28 <= lineBuffer_27;
    end
    if (sel) begin
      lineBuffer_29 <= lineBuffer_28;
    end
    if (sel) begin
      lineBuffer_30 <= lineBuffer_29;
    end
    if (sel) begin
      lineBuffer_31 <= lineBuffer_30;
    end
    if (sel) begin
      lineBuffer_32 <= lineBuffer_31;
    end
    if (sel) begin
      lineBuffer_33 <= lineBuffer_32;
    end
    if (sel) begin
      lineBuffer_34 <= lineBuffer_33;
    end
    if (sel) begin
      lineBuffer_35 <= lineBuffer_34;
    end
    if (sel) begin
      lineBuffer_36 <= lineBuffer_35;
    end
    if (sel) begin
      lineBuffer_37 <= lineBuffer_36;
    end
    if (sel) begin
      lineBuffer_38 <= lineBuffer_37;
    end
    if (sel) begin
      lineBuffer_39 <= lineBuffer_38;
    end
    if (sel) begin
      lineBuffer_40 <= lineBuffer_39;
    end
    if (sel) begin
      lineBuffer_41 <= lineBuffer_40;
    end
    if (sel) begin
      lineBuffer_42 <= lineBuffer_41;
    end
    if (sel) begin
      lineBuffer_43 <= lineBuffer_42;
    end
    if (sel) begin
      lineBuffer_44 <= lineBuffer_43;
    end
    if (sel) begin
      lineBuffer_45 <= lineBuffer_44;
    end
    if (sel) begin
      lineBuffer_46 <= lineBuffer_45;
    end
    if (sel) begin
      lineBuffer_47 <= lineBuffer_46;
    end
    if (sel) begin
      lineBuffer_48 <= lineBuffer_47;
    end
    if (sel) begin
      lineBuffer_49 <= lineBuffer_48;
    end
    if (sel) begin
      lineBuffer_50 <= lineBuffer_49;
    end
    if (sel) begin
      lineBuffer_51 <= lineBuffer_50;
    end
    if (sel) begin
      lineBuffer_52 <= lineBuffer_51;
    end
    if (sel) begin
      lineBuffer_53 <= lineBuffer_52;
    end
    if (sel) begin
      lineBuffer_54 <= lineBuffer_53;
    end
    if (sel) begin
      lineBuffer_55 <= lineBuffer_54;
    end
    if (sel) begin
      lineBuffer_56 <= lineBuffer_55;
    end
    if (sel) begin
      lineBuffer_57 <= lineBuffer_56;
    end
    if (sel) begin
      lineBuffer_58 <= lineBuffer_57;
    end
    if (sel) begin
      lineBuffer_59 <= lineBuffer_58;
    end
    if (sel) begin
      lineBuffer_60 <= lineBuffer_59;
    end
    if (sel) begin
      lineBuffer_61 <= lineBuffer_60;
    end
    if (sel) begin
      lineBuffer_62 <= lineBuffer_61;
    end
    if (sel) begin
      lineBuffer_63 <= lineBuffer_62;
    end
    if (sel) begin
      lineBuffer_64 <= lineBuffer_63;
    end
    if (sel) begin
      lineBuffer_65 <= lineBuffer_64;
    end
    if (sel) begin
      lineBuffer_66 <= lineBuffer_65;
    end
    if (sel) begin
      lineBuffer_67 <= lineBuffer_66;
    end
    if (sel) begin
      lineBuffer_68 <= lineBuffer_67;
    end
    if (sel) begin
      lineBuffer_69 <= lineBuffer_68;
    end
    if (sel) begin
      lineBuffer_70 <= lineBuffer_69;
    end
    if (sel) begin
      lineBuffer_71 <= lineBuffer_70;
    end
    if (sel) begin
      lineBuffer_72 <= lineBuffer_71;
    end
    if (sel) begin
      lineBuffer_73 <= lineBuffer_72;
    end
    if (sel) begin
      lineBuffer_74 <= lineBuffer_73;
    end
    if (sel) begin
      lineBuffer_75 <= lineBuffer_74;
    end
    if (sel) begin
      lineBuffer_76 <= lineBuffer_75;
    end
    if (sel) begin
      lineBuffer_77 <= lineBuffer_76;
    end
    if (sel) begin
      lineBuffer_78 <= lineBuffer_77;
    end
    if (sel) begin
      lineBuffer_79 <= lineBuffer_78;
    end
    if (sel) begin
      lineBuffer_80 <= lineBuffer_79;
    end
    if (sel) begin
      lineBuffer_81 <= lineBuffer_80;
    end
    if (sel) begin
      lineBuffer_82 <= lineBuffer_81;
    end
    if (sel) begin
      lineBuffer_83 <= lineBuffer_82;
    end
    if (sel) begin
      lineBuffer_84 <= lineBuffer_83;
    end
    if (sel) begin
      lineBuffer_85 <= lineBuffer_84;
    end
    if (sel) begin
      lineBuffer_86 <= lineBuffer_85;
    end
    if (sel) begin
      lineBuffer_87 <= lineBuffer_86;
    end
    if (sel) begin
      lineBuffer_88 <= lineBuffer_87;
    end
    if (sel) begin
      lineBuffer_89 <= lineBuffer_88;
    end
    if (sel) begin
      lineBuffer_90 <= lineBuffer_89;
    end
    if (sel) begin
      lineBuffer_91 <= lineBuffer_90;
    end
    if (sel) begin
      lineBuffer_92 <= lineBuffer_91;
    end
    if (sel) begin
      lineBuffer_93 <= lineBuffer_92;
    end
    if (sel) begin
      lineBuffer_94 <= lineBuffer_93;
    end
    if (sel) begin
      lineBuffer_95 <= lineBuffer_94;
    end
    if (sel) begin
      lineBuffer_96 <= lineBuffer_95;
    end
    if (sel) begin
      lineBuffer_97 <= lineBuffer_96;
    end
    if (sel) begin
      lineBuffer_98 <= lineBuffer_97;
    end
    if (sel) begin
      lineBuffer_99 <= lineBuffer_98;
    end
    if (sel) begin
      lineBuffer_100 <= lineBuffer_99;
    end
    if (sel) begin
      lineBuffer_101 <= lineBuffer_100;
    end
    if (sel) begin
      lineBuffer_102 <= lineBuffer_101;
    end
    if (sel) begin
      lineBuffer_103 <= lineBuffer_102;
    end
    if (sel) begin
      lineBuffer_104 <= lineBuffer_103;
    end
    if (sel) begin
      lineBuffer_105 <= lineBuffer_104;
    end
    if (sel) begin
      lineBuffer_106 <= lineBuffer_105;
    end
    if (sel) begin
      lineBuffer_107 <= lineBuffer_106;
    end
    if (sel) begin
      lineBuffer_108 <= lineBuffer_107;
    end
    if (sel) begin
      lineBuffer_109 <= lineBuffer_108;
    end
    if (sel) begin
      lineBuffer_110 <= lineBuffer_109;
    end
    if (sel) begin
      lineBuffer_111 <= lineBuffer_110;
    end
    if (sel) begin
      lineBuffer_112 <= lineBuffer_111;
    end
    if (sel) begin
      lineBuffer_113 <= lineBuffer_112;
    end
    if (sel) begin
      lineBuffer_114 <= lineBuffer_113;
    end
    if (sel) begin
      lineBuffer_115 <= lineBuffer_114;
    end
    if (sel) begin
      lineBuffer_116 <= lineBuffer_115;
    end
    if (sel) begin
      lineBuffer_117 <= lineBuffer_116;
    end
    if (sel) begin
      lineBuffer_118 <= lineBuffer_117;
    end
    if (sel) begin
      lineBuffer_119 <= lineBuffer_118;
    end
    if (sel) begin
      lineBuffer_120 <= lineBuffer_119;
    end
    if (sel) begin
      lineBuffer_121 <= lineBuffer_120;
    end
    if (sel) begin
      lineBuffer_122 <= lineBuffer_121;
    end
    if (sel) begin
      lineBuffer_123 <= lineBuffer_122;
    end
    if (sel) begin
      lineBuffer_124 <= lineBuffer_123;
    end
    if (sel) begin
      lineBuffer_125 <= lineBuffer_124;
    end
    if (sel) begin
      lineBuffer_126 <= lineBuffer_125;
    end
    if (sel) begin
      lineBuffer_127 <= lineBuffer_126;
    end
    if (sel) begin
      lineBuffer_128 <= lineBuffer_127;
    end
    if (sel) begin
      lineBuffer_129 <= lineBuffer_128;
    end
    if (sel) begin
      lineBuffer_130 <= lineBuffer_129;
    end
    if (sel) begin
      lineBuffer_131 <= lineBuffer_130;
    end
    if (sel) begin
      lineBuffer_132 <= lineBuffer_131;
    end
    if (sel) begin
      lineBuffer_133 <= lineBuffer_132;
    end
    if (sel) begin
      lineBuffer_134 <= lineBuffer_133;
    end
    if (sel) begin
      lineBuffer_135 <= lineBuffer_134;
    end
    if (sel) begin
      lineBuffer_136 <= lineBuffer_135;
    end
    if (sel) begin
      lineBuffer_137 <= lineBuffer_136;
    end
    if (sel) begin
      lineBuffer_138 <= lineBuffer_137;
    end
    if (sel) begin
      lineBuffer_139 <= lineBuffer_138;
    end
    if (sel) begin
      lineBuffer_140 <= lineBuffer_139;
    end
    if (sel) begin
      lineBuffer_141 <= lineBuffer_140;
    end
    if (sel) begin
      lineBuffer_142 <= lineBuffer_141;
    end
    if (sel) begin
      lineBuffer_143 <= lineBuffer_142;
    end
    if (sel) begin
      lineBuffer_144 <= lineBuffer_143;
    end
    if (sel) begin
      lineBuffer_145 <= lineBuffer_144;
    end
    if (sel) begin
      lineBuffer_146 <= lineBuffer_145;
    end
    if (sel) begin
      lineBuffer_147 <= lineBuffer_146;
    end
    if (sel) begin
      lineBuffer_148 <= lineBuffer_147;
    end
    if (sel) begin
      lineBuffer_149 <= lineBuffer_148;
    end
    if (sel) begin
      lineBuffer_150 <= lineBuffer_149;
    end
    if (sel) begin
      lineBuffer_151 <= lineBuffer_150;
    end
    if (sel) begin
      lineBuffer_152 <= lineBuffer_151;
    end
    if (sel) begin
      lineBuffer_153 <= lineBuffer_152;
    end
    if (sel) begin
      lineBuffer_154 <= lineBuffer_153;
    end
    if (sel) begin
      lineBuffer_155 <= lineBuffer_154;
    end
    if (sel) begin
      lineBuffer_156 <= lineBuffer_155;
    end
    if (sel) begin
      lineBuffer_157 <= lineBuffer_156;
    end
    if (sel) begin
      lineBuffer_158 <= lineBuffer_157;
    end
    if (sel) begin
      lineBuffer_159 <= lineBuffer_158;
    end
    if (sel) begin
      lineBuffer_160 <= lineBuffer_159;
    end
    if (sel) begin
      lineBuffer_161 <= lineBuffer_160;
    end
    if (sel) begin
      lineBuffer_162 <= lineBuffer_161;
    end
    if (sel) begin
      lineBuffer_163 <= lineBuffer_162;
    end
    if (sel) begin
      lineBuffer_164 <= lineBuffer_163;
    end
    if (sel) begin
      lineBuffer_165 <= lineBuffer_164;
    end
    if (sel) begin
      lineBuffer_166 <= lineBuffer_165;
    end
    if (sel) begin
      lineBuffer_167 <= lineBuffer_166;
    end
    if (sel) begin
      lineBuffer_168 <= lineBuffer_167;
    end
    if (sel) begin
      lineBuffer_169 <= lineBuffer_168;
    end
    if (sel) begin
      lineBuffer_170 <= lineBuffer_169;
    end
    if (sel) begin
      lineBuffer_171 <= lineBuffer_170;
    end
    if (sel) begin
      lineBuffer_172 <= lineBuffer_171;
    end
    if (sel) begin
      lineBuffer_173 <= lineBuffer_172;
    end
    if (sel) begin
      lineBuffer_174 <= lineBuffer_173;
    end
    if (sel) begin
      lineBuffer_175 <= lineBuffer_174;
    end
    if (sel) begin
      lineBuffer_176 <= lineBuffer_175;
    end
    if (sel) begin
      lineBuffer_177 <= lineBuffer_176;
    end
    if (sel) begin
      lineBuffer_178 <= lineBuffer_177;
    end
    if (sel) begin
      lineBuffer_179 <= lineBuffer_178;
    end
    if (sel) begin
      lineBuffer_180 <= lineBuffer_179;
    end
    if (sel) begin
      lineBuffer_181 <= lineBuffer_180;
    end
    if (sel) begin
      lineBuffer_182 <= lineBuffer_181;
    end
    if (sel) begin
      lineBuffer_183 <= lineBuffer_182;
    end
    if (sel) begin
      lineBuffer_184 <= lineBuffer_183;
    end
    if (sel) begin
      lineBuffer_185 <= lineBuffer_184;
    end
    if (sel) begin
      lineBuffer_186 <= lineBuffer_185;
    end
    if (sel) begin
      lineBuffer_187 <= lineBuffer_186;
    end
    if (sel) begin
      lineBuffer_188 <= lineBuffer_187;
    end
    if (sel) begin
      lineBuffer_189 <= lineBuffer_188;
    end
    if (sel) begin
      lineBuffer_190 <= lineBuffer_189;
    end
    if (sel) begin
      lineBuffer_191 <= lineBuffer_190;
    end
    if (sel) begin
      lineBuffer_192 <= lineBuffer_191;
    end
    if (sel) begin
      lineBuffer_193 <= lineBuffer_192;
    end
    if (sel) begin
      lineBuffer_194 <= lineBuffer_193;
    end
    if (sel) begin
      lineBuffer_195 <= lineBuffer_194;
    end
    if (sel) begin
      lineBuffer_196 <= lineBuffer_195;
    end
    if (sel) begin
      lineBuffer_197 <= lineBuffer_196;
    end
    if (sel) begin
      lineBuffer_198 <= lineBuffer_197;
    end
    if (sel) begin
      lineBuffer_199 <= lineBuffer_198;
    end
    if (sel) begin
      lineBuffer_200 <= lineBuffer_199;
    end
    if (sel) begin
      lineBuffer_201 <= lineBuffer_200;
    end
    if (sel) begin
      lineBuffer_202 <= lineBuffer_201;
    end
    if (sel) begin
      lineBuffer_203 <= lineBuffer_202;
    end
    if (sel) begin
      lineBuffer_204 <= lineBuffer_203;
    end
    if (sel) begin
      lineBuffer_205 <= lineBuffer_204;
    end
    if (sel) begin
      lineBuffer_206 <= lineBuffer_205;
    end
    if (sel) begin
      lineBuffer_207 <= lineBuffer_206;
    end
    if (sel) begin
      lineBuffer_208 <= lineBuffer_207;
    end
    if (sel) begin
      lineBuffer_209 <= lineBuffer_208;
    end
    if (sel) begin
      lineBuffer_210 <= lineBuffer_209;
    end
    if (sel) begin
      lineBuffer_211 <= lineBuffer_210;
    end
    if (sel) begin
      lineBuffer_212 <= lineBuffer_211;
    end
    if (sel) begin
      lineBuffer_213 <= lineBuffer_212;
    end
    if (sel) begin
      lineBuffer_214 <= lineBuffer_213;
    end
    if (sel) begin
      lineBuffer_215 <= lineBuffer_214;
    end
    if (sel) begin
      lineBuffer_216 <= lineBuffer_215;
    end
    if (sel) begin
      lineBuffer_217 <= lineBuffer_216;
    end
    if (sel) begin
      lineBuffer_218 <= lineBuffer_217;
    end
    if (sel) begin
      lineBuffer_219 <= lineBuffer_218;
    end
    if (sel) begin
      lineBuffer_220 <= lineBuffer_219;
    end
    if (sel) begin
      lineBuffer_221 <= lineBuffer_220;
    end
    if (sel) begin
      lineBuffer_222 <= lineBuffer_221;
    end
    if (sel) begin
      lineBuffer_223 <= lineBuffer_222;
    end
    if (sel) begin
      lineBuffer_224 <= lineBuffer_223;
    end
    if (sel) begin
      lineBuffer_225 <= lineBuffer_224;
    end
    if (sel) begin
      lineBuffer_226 <= lineBuffer_225;
    end
    if (sel) begin
      lineBuffer_227 <= lineBuffer_226;
    end
    if (sel) begin
      lineBuffer_228 <= lineBuffer_227;
    end
    if (sel) begin
      lineBuffer_229 <= lineBuffer_228;
    end
    if (sel) begin
      lineBuffer_230 <= lineBuffer_229;
    end
    if (sel) begin
      lineBuffer_231 <= lineBuffer_230;
    end
    if (sel) begin
      lineBuffer_232 <= lineBuffer_231;
    end
    if (sel) begin
      lineBuffer_233 <= lineBuffer_232;
    end
    if (sel) begin
      lineBuffer_234 <= lineBuffer_233;
    end
    if (sel) begin
      lineBuffer_235 <= lineBuffer_234;
    end
    if (sel) begin
      lineBuffer_236 <= lineBuffer_235;
    end
    if (sel) begin
      lineBuffer_237 <= lineBuffer_236;
    end
    if (sel) begin
      lineBuffer_238 <= lineBuffer_237;
    end
    if (sel) begin
      lineBuffer_239 <= lineBuffer_238;
    end
    if (sel) begin
      lineBuffer_240 <= lineBuffer_239;
    end
    if (sel) begin
      lineBuffer_241 <= lineBuffer_240;
    end
    if (sel) begin
      lineBuffer_242 <= lineBuffer_241;
    end
    if (sel) begin
      lineBuffer_243 <= lineBuffer_242;
    end
    if (sel) begin
      lineBuffer_244 <= lineBuffer_243;
    end
    if (sel) begin
      lineBuffer_245 <= lineBuffer_244;
    end
    if (sel) begin
      lineBuffer_246 <= lineBuffer_245;
    end
    if (sel) begin
      lineBuffer_247 <= lineBuffer_246;
    end
    if (sel) begin
      lineBuffer_248 <= lineBuffer_247;
    end
    if (sel) begin
      lineBuffer_249 <= lineBuffer_248;
    end
    if (sel) begin
      lineBuffer_250 <= lineBuffer_249;
    end
    if (sel) begin
      lineBuffer_251 <= lineBuffer_250;
    end
    if (sel) begin
      lineBuffer_252 <= lineBuffer_251;
    end
    if (sel) begin
      lineBuffer_253 <= lineBuffer_252;
    end
    if (sel) begin
      lineBuffer_254 <= lineBuffer_253;
    end
    if (sel) begin
      lineBuffer_255 <= lineBuffer_254;
    end
    if (sel) begin
      lineBuffer_256 <= lineBuffer_255;
    end
    if (sel) begin
      lineBuffer_257 <= lineBuffer_256;
    end
    if (sel) begin
      lineBuffer_258 <= lineBuffer_257;
    end
    if (sel) begin
      lineBuffer_259 <= lineBuffer_258;
    end
    if (sel) begin
      lineBuffer_260 <= lineBuffer_259;
    end
    if (sel) begin
      lineBuffer_261 <= lineBuffer_260;
    end
    if (sel) begin
      lineBuffer_262 <= lineBuffer_261;
    end
    if (sel) begin
      lineBuffer_263 <= lineBuffer_262;
    end
    if (sel) begin
      lineBuffer_264 <= lineBuffer_263;
    end
    if (sel) begin
      lineBuffer_265 <= lineBuffer_264;
    end
    if (sel) begin
      lineBuffer_266 <= lineBuffer_265;
    end
    if (sel) begin
      lineBuffer_267 <= lineBuffer_266;
    end
    if (sel) begin
      lineBuffer_268 <= lineBuffer_267;
    end
    if (sel) begin
      lineBuffer_269 <= lineBuffer_268;
    end
    if (sel) begin
      lineBuffer_270 <= lineBuffer_269;
    end
    if (sel) begin
      lineBuffer_271 <= lineBuffer_270;
    end
    if (sel) begin
      lineBuffer_272 <= lineBuffer_271;
    end
    if (sel) begin
      lineBuffer_273 <= lineBuffer_272;
    end
    if (sel) begin
      lineBuffer_274 <= lineBuffer_273;
    end
    if (sel) begin
      lineBuffer_275 <= lineBuffer_274;
    end
    if (sel) begin
      lineBuffer_276 <= lineBuffer_275;
    end
    if (sel) begin
      lineBuffer_277 <= lineBuffer_276;
    end
    if (sel) begin
      lineBuffer_278 <= lineBuffer_277;
    end
    if (sel) begin
      lineBuffer_279 <= lineBuffer_278;
    end
    if (sel) begin
      lineBuffer_280 <= lineBuffer_279;
    end
    if (sel) begin
      lineBuffer_281 <= lineBuffer_280;
    end
    if (sel) begin
      lineBuffer_282 <= lineBuffer_281;
    end
    if (sel) begin
      lineBuffer_283 <= lineBuffer_282;
    end
    if (sel) begin
      lineBuffer_284 <= lineBuffer_283;
    end
    if (sel) begin
      lineBuffer_285 <= lineBuffer_284;
    end
    if (sel) begin
      lineBuffer_286 <= lineBuffer_285;
    end
    if (sel) begin
      lineBuffer_287 <= lineBuffer_286;
    end
    if (sel) begin
      lineBuffer_288 <= lineBuffer_287;
    end
    if (sel) begin
      lineBuffer_289 <= lineBuffer_288;
    end
    if (sel) begin
      lineBuffer_290 <= lineBuffer_289;
    end
    if (sel) begin
      lineBuffer_291 <= lineBuffer_290;
    end
    if (sel) begin
      lineBuffer_292 <= lineBuffer_291;
    end
    if (sel) begin
      lineBuffer_293 <= lineBuffer_292;
    end
    if (sel) begin
      lineBuffer_294 <= lineBuffer_293;
    end
    if (sel) begin
      lineBuffer_295 <= lineBuffer_294;
    end
    if (sel) begin
      lineBuffer_296 <= lineBuffer_295;
    end
    if (sel) begin
      lineBuffer_297 <= lineBuffer_296;
    end
    if (sel) begin
      lineBuffer_298 <= lineBuffer_297;
    end
    if (sel) begin
      lineBuffer_299 <= lineBuffer_298;
    end
    if (sel) begin
      lineBuffer_300 <= lineBuffer_299;
    end
    if (sel) begin
      lineBuffer_301 <= lineBuffer_300;
    end
    if (sel) begin
      lineBuffer_302 <= lineBuffer_301;
    end
    if (sel) begin
      lineBuffer_303 <= lineBuffer_302;
    end
    if (sel) begin
      lineBuffer_304 <= lineBuffer_303;
    end
    if (sel) begin
      lineBuffer_305 <= lineBuffer_304;
    end
    if (sel) begin
      lineBuffer_306 <= lineBuffer_305;
    end
    if (sel) begin
      lineBuffer_307 <= lineBuffer_306;
    end
    if (sel) begin
      lineBuffer_308 <= lineBuffer_307;
    end
    if (sel) begin
      lineBuffer_309 <= lineBuffer_308;
    end
    if (sel) begin
      lineBuffer_310 <= lineBuffer_309;
    end
    if (sel) begin
      lineBuffer_311 <= lineBuffer_310;
    end
    if (sel) begin
      lineBuffer_312 <= lineBuffer_311;
    end
    if (sel) begin
      lineBuffer_313 <= lineBuffer_312;
    end
    if (sel) begin
      lineBuffer_314 <= lineBuffer_313;
    end
    if (sel) begin
      lineBuffer_315 <= lineBuffer_314;
    end
    if (sel) begin
      lineBuffer_316 <= lineBuffer_315;
    end
    if (sel) begin
      lineBuffer_317 <= lineBuffer_316;
    end
    if (sel) begin
      lineBuffer_318 <= lineBuffer_317;
    end
    if (sel) begin
      lineBuffer_319 <= lineBuffer_318;
    end
    if (sel) begin
      lineBuffer_320 <= lineBuffer_319;
    end
    if (sel) begin
      lineBuffer_321 <= lineBuffer_320;
    end
    if (sel) begin
      lineBuffer_322 <= lineBuffer_321;
    end
    if (sel) begin
      lineBuffer_323 <= lineBuffer_322;
    end
    if (sel) begin
      lineBuffer_324 <= lineBuffer_323;
    end
    if (sel) begin
      lineBuffer_325 <= lineBuffer_324;
    end
    if (sel) begin
      lineBuffer_326 <= lineBuffer_325;
    end
    if (sel) begin
      lineBuffer_327 <= lineBuffer_326;
    end
    if (sel) begin
      lineBuffer_328 <= lineBuffer_327;
    end
    if (sel) begin
      lineBuffer_329 <= lineBuffer_328;
    end
    if (sel) begin
      lineBuffer_330 <= lineBuffer_329;
    end
    if (sel) begin
      lineBuffer_331 <= lineBuffer_330;
    end
    if (sel) begin
      lineBuffer_332 <= lineBuffer_331;
    end
    if (sel) begin
      lineBuffer_333 <= lineBuffer_332;
    end
    if (sel) begin
      lineBuffer_334 <= lineBuffer_333;
    end
    if (sel) begin
      lineBuffer_335 <= lineBuffer_334;
    end
    if (sel) begin
      lineBuffer_336 <= lineBuffer_335;
    end
    if (sel) begin
      lineBuffer_337 <= lineBuffer_336;
    end
    if (sel) begin
      lineBuffer_338 <= lineBuffer_337;
    end
    if (sel) begin
      lineBuffer_339 <= lineBuffer_338;
    end
    if (sel) begin
      lineBuffer_340 <= lineBuffer_339;
    end
    if (sel) begin
      lineBuffer_341 <= lineBuffer_340;
    end
    if (sel) begin
      lineBuffer_342 <= lineBuffer_341;
    end
    if (sel) begin
      lineBuffer_343 <= lineBuffer_342;
    end
    if (sel) begin
      lineBuffer_344 <= lineBuffer_343;
    end
    if (sel) begin
      lineBuffer_345 <= lineBuffer_344;
    end
    if (sel) begin
      lineBuffer_346 <= lineBuffer_345;
    end
    if (sel) begin
      lineBuffer_347 <= lineBuffer_346;
    end
    if (sel) begin
      lineBuffer_348 <= lineBuffer_347;
    end
    if (sel) begin
      lineBuffer_349 <= lineBuffer_348;
    end
    if (sel) begin
      lineBuffer_350 <= lineBuffer_349;
    end
    if (sel) begin
      lineBuffer_351 <= lineBuffer_350;
    end
    if (sel) begin
      lineBuffer_352 <= lineBuffer_351;
    end
    if (sel) begin
      lineBuffer_353 <= lineBuffer_352;
    end
    if (sel) begin
      lineBuffer_354 <= lineBuffer_353;
    end
    if (sel) begin
      lineBuffer_355 <= lineBuffer_354;
    end
    if (sel) begin
      lineBuffer_356 <= lineBuffer_355;
    end
    if (sel) begin
      lineBuffer_357 <= lineBuffer_356;
    end
    if (sel) begin
      lineBuffer_358 <= lineBuffer_357;
    end
    if (sel) begin
      lineBuffer_359 <= lineBuffer_358;
    end
    if (sel) begin
      lineBuffer_360 <= lineBuffer_359;
    end
    if (sel) begin
      lineBuffer_361 <= lineBuffer_360;
    end
    if (sel) begin
      lineBuffer_362 <= lineBuffer_361;
    end
    if (sel) begin
      lineBuffer_363 <= lineBuffer_362;
    end
    if (sel) begin
      lineBuffer_364 <= lineBuffer_363;
    end
    if (sel) begin
      lineBuffer_365 <= lineBuffer_364;
    end
    if (sel) begin
      lineBuffer_366 <= lineBuffer_365;
    end
    if (sel) begin
      lineBuffer_367 <= lineBuffer_366;
    end
    if (sel) begin
      lineBuffer_368 <= lineBuffer_367;
    end
    if (sel) begin
      lineBuffer_369 <= lineBuffer_368;
    end
    if (sel) begin
      lineBuffer_370 <= lineBuffer_369;
    end
    if (sel) begin
      lineBuffer_371 <= lineBuffer_370;
    end
    if (sel) begin
      lineBuffer_372 <= lineBuffer_371;
    end
    if (sel) begin
      lineBuffer_373 <= lineBuffer_372;
    end
    if (sel) begin
      lineBuffer_374 <= lineBuffer_373;
    end
    if (sel) begin
      lineBuffer_375 <= lineBuffer_374;
    end
    if (sel) begin
      lineBuffer_376 <= lineBuffer_375;
    end
    if (sel) begin
      lineBuffer_377 <= lineBuffer_376;
    end
    if (sel) begin
      lineBuffer_378 <= lineBuffer_377;
    end
    if (sel) begin
      lineBuffer_379 <= lineBuffer_378;
    end
    if (sel) begin
      lineBuffer_380 <= lineBuffer_379;
    end
    if (sel) begin
      lineBuffer_381 <= lineBuffer_380;
    end
    if (sel) begin
      lineBuffer_382 <= lineBuffer_381;
    end
    if (sel) begin
      lineBuffer_383 <= lineBuffer_382;
    end
    if (sel) begin
      lineBuffer_384 <= lineBuffer_383;
    end
    if (sel) begin
      lineBuffer_385 <= lineBuffer_384;
    end
    if (sel) begin
      lineBuffer_386 <= lineBuffer_385;
    end
    if (sel) begin
      lineBuffer_387 <= lineBuffer_386;
    end
    if (sel) begin
      lineBuffer_388 <= lineBuffer_387;
    end
    if (sel) begin
      lineBuffer_389 <= lineBuffer_388;
    end
    if (sel) begin
      lineBuffer_390 <= lineBuffer_389;
    end
    if (sel) begin
      lineBuffer_391 <= lineBuffer_390;
    end
    if (sel) begin
      lineBuffer_392 <= lineBuffer_391;
    end
    if (sel) begin
      lineBuffer_393 <= lineBuffer_392;
    end
    if (sel) begin
      lineBuffer_394 <= lineBuffer_393;
    end
    if (sel) begin
      lineBuffer_395 <= lineBuffer_394;
    end
    if (sel) begin
      lineBuffer_396 <= lineBuffer_395;
    end
    if (sel) begin
      lineBuffer_397 <= lineBuffer_396;
    end
    if (sel) begin
      lineBuffer_398 <= lineBuffer_397;
    end
    if (sel) begin
      lineBuffer_399 <= lineBuffer_398;
    end
    if (sel) begin
      lineBuffer_400 <= lineBuffer_399;
    end
    if (sel) begin
      lineBuffer_401 <= lineBuffer_400;
    end
    if (sel) begin
      lineBuffer_402 <= lineBuffer_401;
    end
    if (sel) begin
      lineBuffer_403 <= lineBuffer_402;
    end
    if (sel) begin
      lineBuffer_404 <= lineBuffer_403;
    end
    if (sel) begin
      lineBuffer_405 <= lineBuffer_404;
    end
    if (sel) begin
      lineBuffer_406 <= lineBuffer_405;
    end
    if (sel) begin
      lineBuffer_407 <= lineBuffer_406;
    end
    if (sel) begin
      lineBuffer_408 <= lineBuffer_407;
    end
    if (sel) begin
      lineBuffer_409 <= lineBuffer_408;
    end
    if (sel) begin
      lineBuffer_410 <= lineBuffer_409;
    end
    if (sel) begin
      lineBuffer_411 <= lineBuffer_410;
    end
    if (sel) begin
      lineBuffer_412 <= lineBuffer_411;
    end
    if (sel) begin
      lineBuffer_413 <= lineBuffer_412;
    end
    if (sel) begin
      lineBuffer_414 <= lineBuffer_413;
    end
    if (sel) begin
      lineBuffer_415 <= lineBuffer_414;
    end
    if (sel) begin
      lineBuffer_416 <= lineBuffer_415;
    end
    if (sel) begin
      lineBuffer_417 <= lineBuffer_416;
    end
    if (sel) begin
      lineBuffer_418 <= lineBuffer_417;
    end
    if (sel) begin
      lineBuffer_419 <= lineBuffer_418;
    end
    if (sel) begin
      lineBuffer_420 <= lineBuffer_419;
    end
    if (sel) begin
      lineBuffer_421 <= lineBuffer_420;
    end
    if (sel) begin
      lineBuffer_422 <= lineBuffer_421;
    end
    if (sel) begin
      lineBuffer_423 <= lineBuffer_422;
    end
    if (sel) begin
      lineBuffer_424 <= lineBuffer_423;
    end
    if (sel) begin
      lineBuffer_425 <= lineBuffer_424;
    end
    if (sel) begin
      lineBuffer_426 <= lineBuffer_425;
    end
    if (sel) begin
      lineBuffer_427 <= lineBuffer_426;
    end
    if (sel) begin
      lineBuffer_428 <= lineBuffer_427;
    end
    if (sel) begin
      lineBuffer_429 <= lineBuffer_428;
    end
    if (sel) begin
      lineBuffer_430 <= lineBuffer_429;
    end
    if (sel) begin
      lineBuffer_431 <= lineBuffer_430;
    end
    if (sel) begin
      lineBuffer_432 <= lineBuffer_431;
    end
    if (sel) begin
      lineBuffer_433 <= lineBuffer_432;
    end
    if (sel) begin
      lineBuffer_434 <= lineBuffer_433;
    end
    if (sel) begin
      lineBuffer_435 <= lineBuffer_434;
    end
    if (sel) begin
      lineBuffer_436 <= lineBuffer_435;
    end
    if (sel) begin
      lineBuffer_437 <= lineBuffer_436;
    end
    if (sel) begin
      lineBuffer_438 <= lineBuffer_437;
    end
    if (sel) begin
      lineBuffer_439 <= lineBuffer_438;
    end
    if (sel) begin
      lineBuffer_440 <= lineBuffer_439;
    end
    if (sel) begin
      lineBuffer_441 <= lineBuffer_440;
    end
    if (sel) begin
      lineBuffer_442 <= lineBuffer_441;
    end
    if (sel) begin
      lineBuffer_443 <= lineBuffer_442;
    end
    if (sel) begin
      lineBuffer_444 <= lineBuffer_443;
    end
    if (sel) begin
      lineBuffer_445 <= lineBuffer_444;
    end
    if (sel) begin
      lineBuffer_446 <= lineBuffer_445;
    end
    if (sel) begin
      lineBuffer_447 <= lineBuffer_446;
    end
    if (sel) begin
      lineBuffer_448 <= lineBuffer_447;
    end
    if (sel) begin
      lineBuffer_449 <= lineBuffer_448;
    end
    if (sel) begin
      lineBuffer_450 <= lineBuffer_449;
    end
    if (sel) begin
      lineBuffer_451 <= lineBuffer_450;
    end
    if (sel) begin
      lineBuffer_452 <= lineBuffer_451;
    end
    if (sel) begin
      lineBuffer_453 <= lineBuffer_452;
    end
    if (sel) begin
      lineBuffer_454 <= lineBuffer_453;
    end
    if (sel) begin
      lineBuffer_455 <= lineBuffer_454;
    end
    if (sel) begin
      lineBuffer_456 <= lineBuffer_455;
    end
    if (sel) begin
      lineBuffer_457 <= lineBuffer_456;
    end
    if (sel) begin
      lineBuffer_458 <= lineBuffer_457;
    end
    if (sel) begin
      lineBuffer_459 <= lineBuffer_458;
    end
    if (sel) begin
      lineBuffer_460 <= lineBuffer_459;
    end
    if (sel) begin
      lineBuffer_461 <= lineBuffer_460;
    end
    if (sel) begin
      lineBuffer_462 <= lineBuffer_461;
    end
    if (sel) begin
      lineBuffer_463 <= lineBuffer_462;
    end
    if (sel) begin
      lineBuffer_464 <= lineBuffer_463;
    end
    if (sel) begin
      lineBuffer_465 <= lineBuffer_464;
    end
    if (sel) begin
      lineBuffer_466 <= lineBuffer_465;
    end
    if (sel) begin
      lineBuffer_467 <= lineBuffer_466;
    end
    if (sel) begin
      lineBuffer_468 <= lineBuffer_467;
    end
    if (sel) begin
      lineBuffer_469 <= lineBuffer_468;
    end
    if (sel) begin
      lineBuffer_470 <= lineBuffer_469;
    end
    if (sel) begin
      lineBuffer_471 <= lineBuffer_470;
    end
    if (sel) begin
      lineBuffer_472 <= lineBuffer_471;
    end
    if (sel) begin
      lineBuffer_473 <= lineBuffer_472;
    end
    if (sel) begin
      lineBuffer_474 <= lineBuffer_473;
    end
    if (sel) begin
      lineBuffer_475 <= lineBuffer_474;
    end
    if (sel) begin
      lineBuffer_476 <= lineBuffer_475;
    end
    if (sel) begin
      lineBuffer_477 <= lineBuffer_476;
    end
    if (sel) begin
      lineBuffer_478 <= lineBuffer_477;
    end
    if (sel) begin
      lineBuffer_479 <= lineBuffer_478;
    end
    if (sel) begin
      lineBuffer_480 <= lineBuffer_479;
    end
    if (sel) begin
      lineBuffer_481 <= lineBuffer_480;
    end
    if (sel) begin
      lineBuffer_482 <= lineBuffer_481;
    end
    if (sel) begin
      lineBuffer_483 <= lineBuffer_482;
    end
    if (sel) begin
      lineBuffer_484 <= lineBuffer_483;
    end
    if (sel) begin
      lineBuffer_485 <= lineBuffer_484;
    end
    if (sel) begin
      lineBuffer_486 <= lineBuffer_485;
    end
    if (sel) begin
      lineBuffer_487 <= lineBuffer_486;
    end
    if (sel) begin
      lineBuffer_488 <= lineBuffer_487;
    end
    if (sel) begin
      lineBuffer_489 <= lineBuffer_488;
    end
    if (sel) begin
      lineBuffer_490 <= lineBuffer_489;
    end
    if (sel) begin
      lineBuffer_491 <= lineBuffer_490;
    end
    if (sel) begin
      lineBuffer_492 <= lineBuffer_491;
    end
    if (sel) begin
      lineBuffer_493 <= lineBuffer_492;
    end
    if (sel) begin
      lineBuffer_494 <= lineBuffer_493;
    end
    if (sel) begin
      lineBuffer_495 <= lineBuffer_494;
    end
    if (sel) begin
      lineBuffer_496 <= lineBuffer_495;
    end
    if (sel) begin
      lineBuffer_497 <= lineBuffer_496;
    end
    if (sel) begin
      lineBuffer_498 <= lineBuffer_497;
    end
    if (sel) begin
      lineBuffer_499 <= lineBuffer_498;
    end
    if (sel) begin
      lineBuffer_500 <= lineBuffer_499;
    end
    if (sel) begin
      lineBuffer_501 <= lineBuffer_500;
    end
    if (sel) begin
      lineBuffer_502 <= lineBuffer_501;
    end
    if (sel) begin
      lineBuffer_503 <= lineBuffer_502;
    end
    if (sel) begin
      lineBuffer_504 <= lineBuffer_503;
    end
    if (sel) begin
      lineBuffer_505 <= lineBuffer_504;
    end
    if (sel) begin
      lineBuffer_506 <= lineBuffer_505;
    end
    if (sel) begin
      lineBuffer_507 <= lineBuffer_506;
    end
    if (sel) begin
      lineBuffer_508 <= lineBuffer_507;
    end
    if (sel) begin
      lineBuffer_509 <= lineBuffer_508;
    end
    if (sel) begin
      lineBuffer_510 <= lineBuffer_509;
    end
    if (sel) begin
      lineBuffer_511 <= lineBuffer_510;
    end
    if (sel) begin
      lineBuffer_512 <= lineBuffer_511;
    end
    if (sel) begin
      lineBuffer_513 <= lineBuffer_512;
    end
    if (sel) begin
      lineBuffer_514 <= lineBuffer_513;
    end
    if (sel) begin
      lineBuffer_515 <= lineBuffer_514;
    end
    if (sel) begin
      lineBuffer_516 <= lineBuffer_515;
    end
    if (sel) begin
      lineBuffer_517 <= lineBuffer_516;
    end
    if (sel) begin
      lineBuffer_518 <= lineBuffer_517;
    end
    if (sel) begin
      lineBuffer_519 <= lineBuffer_518;
    end
    if (sel) begin
      lineBuffer_520 <= lineBuffer_519;
    end
    if (sel) begin
      lineBuffer_521 <= lineBuffer_520;
    end
    if (sel) begin
      lineBuffer_522 <= lineBuffer_521;
    end
    if (sel) begin
      lineBuffer_523 <= lineBuffer_522;
    end
    if (sel) begin
      lineBuffer_524 <= lineBuffer_523;
    end
    if (sel) begin
      lineBuffer_525 <= lineBuffer_524;
    end
    if (sel) begin
      lineBuffer_526 <= lineBuffer_525;
    end
    if (sel) begin
      lineBuffer_527 <= lineBuffer_526;
    end
    if (sel) begin
      lineBuffer_528 <= lineBuffer_527;
    end
    if (sel) begin
      lineBuffer_529 <= lineBuffer_528;
    end
    if (sel) begin
      lineBuffer_530 <= lineBuffer_529;
    end
    if (sel) begin
      lineBuffer_531 <= lineBuffer_530;
    end
    if (sel) begin
      lineBuffer_532 <= lineBuffer_531;
    end
    if (sel) begin
      lineBuffer_533 <= lineBuffer_532;
    end
    if (sel) begin
      lineBuffer_534 <= lineBuffer_533;
    end
    if (sel) begin
      lineBuffer_535 <= lineBuffer_534;
    end
    if (sel) begin
      lineBuffer_536 <= lineBuffer_535;
    end
    if (sel) begin
      lineBuffer_537 <= lineBuffer_536;
    end
    if (sel) begin
      lineBuffer_538 <= lineBuffer_537;
    end
    if (sel) begin
      lineBuffer_539 <= lineBuffer_538;
    end
    if (sel) begin
      lineBuffer_540 <= lineBuffer_539;
    end
    if (sel) begin
      lineBuffer_541 <= lineBuffer_540;
    end
    if (sel) begin
      lineBuffer_542 <= lineBuffer_541;
    end
    if (sel) begin
      lineBuffer_543 <= lineBuffer_542;
    end
    if (sel) begin
      lineBuffer_544 <= lineBuffer_543;
    end
    if (sel) begin
      lineBuffer_545 <= lineBuffer_544;
    end
    if (sel) begin
      lineBuffer_546 <= lineBuffer_545;
    end
    if (sel) begin
      lineBuffer_547 <= lineBuffer_546;
    end
    if (sel) begin
      lineBuffer_548 <= lineBuffer_547;
    end
    if (sel) begin
      lineBuffer_549 <= lineBuffer_548;
    end
    if (sel) begin
      lineBuffer_550 <= lineBuffer_549;
    end
    if (sel) begin
      lineBuffer_551 <= lineBuffer_550;
    end
    if (sel) begin
      lineBuffer_552 <= lineBuffer_551;
    end
    if (sel) begin
      lineBuffer_553 <= lineBuffer_552;
    end
    if (sel) begin
      lineBuffer_554 <= lineBuffer_553;
    end
    if (sel) begin
      lineBuffer_555 <= lineBuffer_554;
    end
    if (sel) begin
      lineBuffer_556 <= lineBuffer_555;
    end
    if (sel) begin
      lineBuffer_557 <= lineBuffer_556;
    end
    if (sel) begin
      lineBuffer_558 <= lineBuffer_557;
    end
    if (sel) begin
      lineBuffer_559 <= lineBuffer_558;
    end
    if (sel) begin
      lineBuffer_560 <= lineBuffer_559;
    end
    if (sel) begin
      lineBuffer_561 <= lineBuffer_560;
    end
    if (sel) begin
      lineBuffer_562 <= lineBuffer_561;
    end
    if (sel) begin
      lineBuffer_563 <= lineBuffer_562;
    end
    if (sel) begin
      lineBuffer_564 <= lineBuffer_563;
    end
    if (sel) begin
      lineBuffer_565 <= lineBuffer_564;
    end
    if (sel) begin
      lineBuffer_566 <= lineBuffer_565;
    end
    if (sel) begin
      lineBuffer_567 <= lineBuffer_566;
    end
    if (sel) begin
      lineBuffer_568 <= lineBuffer_567;
    end
    if (sel) begin
      lineBuffer_569 <= lineBuffer_568;
    end
    if (sel) begin
      lineBuffer_570 <= lineBuffer_569;
    end
    if (sel) begin
      lineBuffer_571 <= lineBuffer_570;
    end
    if (sel) begin
      lineBuffer_572 <= lineBuffer_571;
    end
    if (sel) begin
      lineBuffer_573 <= lineBuffer_572;
    end
    if (sel) begin
      lineBuffer_574 <= lineBuffer_573;
    end
    if (sel) begin
      lineBuffer_575 <= lineBuffer_574;
    end
    if (sel) begin
      lineBuffer_576 <= lineBuffer_575;
    end
    if (sel) begin
      lineBuffer_577 <= lineBuffer_576;
    end
    if (sel) begin
      lineBuffer_578 <= lineBuffer_577;
    end
    if (sel) begin
      lineBuffer_579 <= lineBuffer_578;
    end
    if (sel) begin
      lineBuffer_580 <= lineBuffer_579;
    end
    if (sel) begin
      lineBuffer_581 <= lineBuffer_580;
    end
    if (sel) begin
      lineBuffer_582 <= lineBuffer_581;
    end
    if (sel) begin
      lineBuffer_583 <= lineBuffer_582;
    end
    if (sel) begin
      lineBuffer_584 <= lineBuffer_583;
    end
    if (sel) begin
      lineBuffer_585 <= lineBuffer_584;
    end
    if (sel) begin
      lineBuffer_586 <= lineBuffer_585;
    end
    if (sel) begin
      lineBuffer_587 <= lineBuffer_586;
    end
    if (sel) begin
      lineBuffer_588 <= lineBuffer_587;
    end
    if (sel) begin
      lineBuffer_589 <= lineBuffer_588;
    end
    if (sel) begin
      lineBuffer_590 <= lineBuffer_589;
    end
    if (sel) begin
      lineBuffer_591 <= lineBuffer_590;
    end
    if (sel) begin
      lineBuffer_592 <= lineBuffer_591;
    end
    if (sel) begin
      lineBuffer_593 <= lineBuffer_592;
    end
    if (sel) begin
      lineBuffer_594 <= lineBuffer_593;
    end
    if (sel) begin
      lineBuffer_595 <= lineBuffer_594;
    end
    if (sel) begin
      lineBuffer_596 <= lineBuffer_595;
    end
    if (sel) begin
      lineBuffer_597 <= lineBuffer_596;
    end
    if (sel) begin
      lineBuffer_598 <= lineBuffer_597;
    end
    if (sel) begin
      lineBuffer_599 <= lineBuffer_598;
    end
    if (sel) begin
      lineBuffer_600 <= lineBuffer_599;
    end
    if (sel) begin
      lineBuffer_601 <= lineBuffer_600;
    end
    if (sel) begin
      lineBuffer_602 <= lineBuffer_601;
    end
    if (sel) begin
      lineBuffer_603 <= lineBuffer_602;
    end
    if (sel) begin
      lineBuffer_604 <= lineBuffer_603;
    end
    if (sel) begin
      lineBuffer_605 <= lineBuffer_604;
    end
    if (sel) begin
      lineBuffer_606 <= lineBuffer_605;
    end
    if (sel) begin
      lineBuffer_607 <= lineBuffer_606;
    end
    if (sel) begin
      lineBuffer_608 <= lineBuffer_607;
    end
    if (sel) begin
      lineBuffer_609 <= lineBuffer_608;
    end
    if (sel) begin
      lineBuffer_610 <= lineBuffer_609;
    end
    if (sel) begin
      lineBuffer_611 <= lineBuffer_610;
    end
    if (sel) begin
      lineBuffer_612 <= lineBuffer_611;
    end
    if (sel) begin
      lineBuffer_613 <= lineBuffer_612;
    end
    if (sel) begin
      lineBuffer_614 <= lineBuffer_613;
    end
    if (sel) begin
      lineBuffer_615 <= lineBuffer_614;
    end
    if (sel) begin
      lineBuffer_616 <= lineBuffer_615;
    end
    if (sel) begin
      lineBuffer_617 <= lineBuffer_616;
    end
    if (sel) begin
      lineBuffer_618 <= lineBuffer_617;
    end
    if (sel) begin
      lineBuffer_619 <= lineBuffer_618;
    end
    if (sel) begin
      lineBuffer_620 <= lineBuffer_619;
    end
    if (sel) begin
      lineBuffer_621 <= lineBuffer_620;
    end
    if (sel) begin
      lineBuffer_622 <= lineBuffer_621;
    end
    if (sel) begin
      lineBuffer_623 <= lineBuffer_622;
    end
    if (sel) begin
      lineBuffer_624 <= lineBuffer_623;
    end
    if (sel) begin
      lineBuffer_625 <= lineBuffer_624;
    end
    if (sel) begin
      lineBuffer_626 <= lineBuffer_625;
    end
    if (sel) begin
      lineBuffer_627 <= lineBuffer_626;
    end
    if (sel) begin
      lineBuffer_628 <= lineBuffer_627;
    end
    if (sel) begin
      lineBuffer_629 <= lineBuffer_628;
    end
    if (sel) begin
      lineBuffer_630 <= lineBuffer_629;
    end
    if (sel) begin
      lineBuffer_631 <= lineBuffer_630;
    end
    if (sel) begin
      lineBuffer_632 <= lineBuffer_631;
    end
    if (sel) begin
      lineBuffer_633 <= lineBuffer_632;
    end
    if (sel) begin
      lineBuffer_634 <= lineBuffer_633;
    end
    if (sel) begin
      lineBuffer_635 <= lineBuffer_634;
    end
    if (sel) begin
      lineBuffer_636 <= lineBuffer_635;
    end
    if (sel) begin
      lineBuffer_637 <= lineBuffer_636;
    end
    if (sel) begin
      lineBuffer_638 <= lineBuffer_637;
    end
    if (sel) begin
      lineBuffer_639 <= lineBuffer_638;
    end
    if (sel) begin
      lineBuffer_640 <= lineBuffer_639;
    end
    if (sel) begin
      lineBuffer_641 <= lineBuffer_640;
    end
    if (sel) begin
      lineBuffer_642 <= lineBuffer_641;
    end
    if (sel) begin
      lineBuffer_643 <= lineBuffer_642;
    end
    if (sel) begin
      lineBuffer_644 <= lineBuffer_643;
    end
    if (sel) begin
      lineBuffer_645 <= lineBuffer_644;
    end
    if (sel) begin
      lineBuffer_646 <= lineBuffer_645;
    end
    if (sel) begin
      lineBuffer_647 <= lineBuffer_646;
    end
    if (sel) begin
      lineBuffer_648 <= lineBuffer_647;
    end
    if (sel) begin
      lineBuffer_649 <= lineBuffer_648;
    end
    if (sel) begin
      lineBuffer_650 <= lineBuffer_649;
    end
    if (sel) begin
      lineBuffer_651 <= lineBuffer_650;
    end
    if (sel) begin
      lineBuffer_652 <= lineBuffer_651;
    end
    if (sel) begin
      lineBuffer_653 <= lineBuffer_652;
    end
    if (sel) begin
      lineBuffer_654 <= lineBuffer_653;
    end
    if (sel) begin
      lineBuffer_655 <= lineBuffer_654;
    end
    if (sel) begin
      lineBuffer_656 <= lineBuffer_655;
    end
    if (sel) begin
      lineBuffer_657 <= lineBuffer_656;
    end
    if (sel) begin
      lineBuffer_658 <= lineBuffer_657;
    end
    if (sel) begin
      lineBuffer_659 <= lineBuffer_658;
    end
    if (sel) begin
      lineBuffer_660 <= lineBuffer_659;
    end
    if (sel) begin
      lineBuffer_661 <= lineBuffer_660;
    end
    if (sel) begin
      lineBuffer_662 <= lineBuffer_661;
    end
    if (sel) begin
      lineBuffer_663 <= lineBuffer_662;
    end
    if (sel) begin
      lineBuffer_664 <= lineBuffer_663;
    end
    if (sel) begin
      lineBuffer_665 <= lineBuffer_664;
    end
    if (sel) begin
      lineBuffer_666 <= lineBuffer_665;
    end
    if (sel) begin
      lineBuffer_667 <= lineBuffer_666;
    end
    if (sel) begin
      lineBuffer_668 <= lineBuffer_667;
    end
    if (sel) begin
      lineBuffer_669 <= lineBuffer_668;
    end
    if (sel) begin
      lineBuffer_670 <= lineBuffer_669;
    end
    if (sel) begin
      lineBuffer_671 <= lineBuffer_670;
    end
    if (sel) begin
      lineBuffer_672 <= lineBuffer_671;
    end
    if (sel) begin
      lineBuffer_673 <= lineBuffer_672;
    end
    if (sel) begin
      lineBuffer_674 <= lineBuffer_673;
    end
    if (sel) begin
      lineBuffer_675 <= lineBuffer_674;
    end
    if (sel) begin
      lineBuffer_676 <= lineBuffer_675;
    end
    if (sel) begin
      lineBuffer_677 <= lineBuffer_676;
    end
    if (sel) begin
      lineBuffer_678 <= lineBuffer_677;
    end
    if (sel) begin
      lineBuffer_679 <= lineBuffer_678;
    end
    if (sel) begin
      lineBuffer_680 <= lineBuffer_679;
    end
    if (sel) begin
      lineBuffer_681 <= lineBuffer_680;
    end
    if (sel) begin
      lineBuffer_682 <= lineBuffer_681;
    end
    if (sel) begin
      lineBuffer_683 <= lineBuffer_682;
    end
    if (sel) begin
      lineBuffer_684 <= lineBuffer_683;
    end
    if (sel) begin
      lineBuffer_685 <= lineBuffer_684;
    end
    if (sel) begin
      lineBuffer_686 <= lineBuffer_685;
    end
    if (sel) begin
      lineBuffer_687 <= lineBuffer_686;
    end
    if (sel) begin
      lineBuffer_688 <= lineBuffer_687;
    end
    if (sel) begin
      lineBuffer_689 <= lineBuffer_688;
    end
    if (sel) begin
      lineBuffer_690 <= lineBuffer_689;
    end
    if (sel) begin
      lineBuffer_691 <= lineBuffer_690;
    end
    if (sel) begin
      lineBuffer_692 <= lineBuffer_691;
    end
    if (sel) begin
      lineBuffer_693 <= lineBuffer_692;
    end
    if (sel) begin
      lineBuffer_694 <= lineBuffer_693;
    end
    if (sel) begin
      lineBuffer_695 <= lineBuffer_694;
    end
    if (sel) begin
      lineBuffer_696 <= lineBuffer_695;
    end
    if (sel) begin
      lineBuffer_697 <= lineBuffer_696;
    end
    if (sel) begin
      lineBuffer_698 <= lineBuffer_697;
    end
    if (sel) begin
      lineBuffer_699 <= lineBuffer_698;
    end
    if (sel) begin
      lineBuffer_700 <= lineBuffer_699;
    end
    if (sel) begin
      lineBuffer_701 <= lineBuffer_700;
    end
    if (sel) begin
      lineBuffer_702 <= lineBuffer_701;
    end
    if (sel) begin
      lineBuffer_703 <= lineBuffer_702;
    end
    if (sel) begin
      lineBuffer_704 <= lineBuffer_703;
    end
    if (sel) begin
      lineBuffer_705 <= lineBuffer_704;
    end
    if (sel) begin
      lineBuffer_706 <= lineBuffer_705;
    end
    if (sel) begin
      lineBuffer_707 <= lineBuffer_706;
    end
    if (sel) begin
      lineBuffer_708 <= lineBuffer_707;
    end
    if (sel) begin
      lineBuffer_709 <= lineBuffer_708;
    end
    if (sel) begin
      lineBuffer_710 <= lineBuffer_709;
    end
    if (sel) begin
      lineBuffer_711 <= lineBuffer_710;
    end
    if (sel) begin
      lineBuffer_712 <= lineBuffer_711;
    end
    if (sel) begin
      lineBuffer_713 <= lineBuffer_712;
    end
    if (sel) begin
      lineBuffer_714 <= lineBuffer_713;
    end
    if (sel) begin
      lineBuffer_715 <= lineBuffer_714;
    end
    if (sel) begin
      lineBuffer_716 <= lineBuffer_715;
    end
    if (sel) begin
      lineBuffer_717 <= lineBuffer_716;
    end
    if (sel) begin
      lineBuffer_718 <= lineBuffer_717;
    end
    if (sel) begin
      lineBuffer_719 <= lineBuffer_718;
    end
    if (sel) begin
      lineBuffer_720 <= lineBuffer_719;
    end
    if (sel) begin
      lineBuffer_721 <= lineBuffer_720;
    end
    if (sel) begin
      lineBuffer_722 <= lineBuffer_721;
    end
    if (sel) begin
      lineBuffer_723 <= lineBuffer_722;
    end
    if (sel) begin
      lineBuffer_724 <= lineBuffer_723;
    end
    if (sel) begin
      lineBuffer_725 <= lineBuffer_724;
    end
    if (sel) begin
      lineBuffer_726 <= lineBuffer_725;
    end
    if (sel) begin
      lineBuffer_727 <= lineBuffer_726;
    end
    if (sel) begin
      lineBuffer_728 <= lineBuffer_727;
    end
    if (sel) begin
      lineBuffer_729 <= lineBuffer_728;
    end
    if (sel) begin
      lineBuffer_730 <= lineBuffer_729;
    end
    if (sel) begin
      lineBuffer_731 <= lineBuffer_730;
    end
    if (sel) begin
      lineBuffer_732 <= lineBuffer_731;
    end
    if (sel) begin
      lineBuffer_733 <= lineBuffer_732;
    end
    if (sel) begin
      lineBuffer_734 <= lineBuffer_733;
    end
    if (sel) begin
      lineBuffer_735 <= lineBuffer_734;
    end
    if (sel) begin
      lineBuffer_736 <= lineBuffer_735;
    end
    if (sel) begin
      lineBuffer_737 <= lineBuffer_736;
    end
    if (sel) begin
      lineBuffer_738 <= lineBuffer_737;
    end
    if (sel) begin
      lineBuffer_739 <= lineBuffer_738;
    end
    if (sel) begin
      lineBuffer_740 <= lineBuffer_739;
    end
    if (sel) begin
      lineBuffer_741 <= lineBuffer_740;
    end
    if (sel) begin
      lineBuffer_742 <= lineBuffer_741;
    end
    if (sel) begin
      lineBuffer_743 <= lineBuffer_742;
    end
    if (sel) begin
      lineBuffer_744 <= lineBuffer_743;
    end
    if (sel) begin
      lineBuffer_745 <= lineBuffer_744;
    end
    if (sel) begin
      lineBuffer_746 <= lineBuffer_745;
    end
    if (sel) begin
      lineBuffer_747 <= lineBuffer_746;
    end
    if (sel) begin
      lineBuffer_748 <= lineBuffer_747;
    end
    if (sel) begin
      lineBuffer_749 <= lineBuffer_748;
    end
    if (sel) begin
      lineBuffer_750 <= lineBuffer_749;
    end
    if (sel) begin
      lineBuffer_751 <= lineBuffer_750;
    end
    if (sel) begin
      lineBuffer_752 <= lineBuffer_751;
    end
    if (sel) begin
      lineBuffer_753 <= lineBuffer_752;
    end
    if (sel) begin
      lineBuffer_754 <= lineBuffer_753;
    end
    if (sel) begin
      lineBuffer_755 <= lineBuffer_754;
    end
    if (sel) begin
      lineBuffer_756 <= lineBuffer_755;
    end
    if (sel) begin
      lineBuffer_757 <= lineBuffer_756;
    end
    if (sel) begin
      lineBuffer_758 <= lineBuffer_757;
    end
    if (sel) begin
      lineBuffer_759 <= lineBuffer_758;
    end
    if (sel) begin
      lineBuffer_760 <= lineBuffer_759;
    end
    if (sel) begin
      lineBuffer_761 <= lineBuffer_760;
    end
    if (sel) begin
      lineBuffer_762 <= lineBuffer_761;
    end
    if (sel) begin
      lineBuffer_763 <= lineBuffer_762;
    end
    if (sel) begin
      lineBuffer_764 <= lineBuffer_763;
    end
    if (sel) begin
      lineBuffer_765 <= lineBuffer_764;
    end
    if (sel) begin
      lineBuffer_766 <= lineBuffer_765;
    end
    if (sel) begin
      lineBuffer_767 <= lineBuffer_766;
    end
    if (sel) begin
      windowBuffer_0 <= windowBuffer_1;
    end
    if (sel) begin
      windowBuffer_1 <= windowBuffer_2;
    end
    if (sel) begin
      windowBuffer_2 <= lineBuffer_255;
    end
    if (sel) begin
      windowBuffer_3 <= windowBuffer_4;
    end
    if (sel) begin
      windowBuffer_4 <= windowBuffer_5;
    end
    if (sel) begin
      windowBuffer_5 <= lineBuffer_511;
    end
    if (sel) begin
      windowBuffer_6 <= windowBuffer_7;
    end
    if (sel) begin
      windowBuffer_7 <= windowBuffer_8;
    end
    if (sel) begin
      windowBuffer_8 <= lineBuffer_767;
    end
  end
endmodule
module Gray2RGBFilter(
  input         clock,
  input         reset,
  output        io_enq_ready,
  input         io_enq_valid,
  input  [23:0] io_enq_bits,
  input         io_enq_user,
  input         io_enq_last,
  input         io_deq_ready,
  output        io_deq_valid,
  output [23:0] io_deq_bits,
  output        io_deq_user,
  output        io_deq_last
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
`endif // RANDOMIZE_REG_INIT
  reg [1:0] stateReg; // @[ChiselImProc.scala 62:28]
  reg [23:0] dataReg; // @[ChiselImProc.scala 64:23]
  reg [23:0] shadowReg; // @[ChiselImProc.scala 66:25]
  reg  userReg; // @[ChiselImProc.scala 67:23]
  reg  shadowUserReg; // @[ChiselImProc.scala 68:29]
  reg  lastReg; // @[ChiselImProc.scala 69:23]
  reg  shadowLastReg; // @[ChiselImProc.scala 70:29]
  wire  _T = 2'h0 == stateReg; // @[Conditional.scala 37:30]
  wire  _T_1 = 2'h1 == stateReg; // @[Conditional.scala 37:30]
  wire  _T_2 = ~io_enq_valid; // @[ChiselImProc.scala 84:39]
  wire  _T_3 = io_deq_ready & _T_2; // @[ChiselImProc.scala 84:36]
  wire  _T_4 = io_deq_ready & io_enq_valid; // @[ChiselImProc.scala 87:42]
  wire  _T_5 = ~io_deq_ready; // @[ChiselImProc.scala 92:29]
  wire  _T_6 = _T_5 & io_enq_valid; // @[ChiselImProc.scala 92:43]
  wire  _T_7 = 2'h2 == stateReg; // @[Conditional.scala 37:30]
  wire  _T_8 = 2'h3 == stateReg; // @[Conditional.scala 37:30]
  wire  _T_9 = stateReg == 2'h0; // @[ChiselImProc.scala 116:35]
  wire  _T_10 = stateReg == 2'h1; // @[ChiselImProc.scala 116:57]
  wire  _T_11 = _T_9 | _T_10; // @[ChiselImProc.scala 116:45]
  wire  _T_12 = stateReg == 2'h3; // @[ChiselImProc.scala 116:77]
  wire  _T_15 = stateReg == 2'h2; // @[ChiselImProc.scala 117:55]
  wire [39:0] _GEN_44 = {dataReg, 16'h0}; // @[ChiselImProc.scala 201:28]
  wire [54:0] _T_17 = {{15'd0}, _GEN_44}; // @[ChiselImProc.scala 201:28]
  wire [31:0] _GEN_45 = {dataReg, 8'h0}; // @[ChiselImProc.scala 201:46]
  wire [38:0] _T_18 = {{7'd0}, _GEN_45}; // @[ChiselImProc.scala 201:46]
  wire [54:0] _GEN_46 = {{16'd0}, _T_18}; // @[ChiselImProc.scala 201:36]
  wire [54:0] _T_19 = _T_17 | _GEN_46; // @[ChiselImProc.scala 201:36]
  wire [54:0] _GEN_47 = {{31'd0}, dataReg}; // @[ChiselImProc.scala 201:53]
  wire [54:0] _T_20 = _T_19 | _GEN_47; // @[ChiselImProc.scala 201:53]
  assign io_enq_ready = _T_11 | _T_12; // @[ChiselImProc.scala 116:22]
  assign io_deq_valid = _T_10 | _T_15; // @[ChiselImProc.scala 117:22]
  assign io_deq_bits = _T_20[23:0]; // @[ChiselImProc.scala 201:17]
  assign io_deq_user = userReg; // @[ChiselImProc.scala 144:17 ChiselImProc.scala 114:21]
  assign io_deq_last = lastReg; // @[ChiselImProc.scala 143:17 ChiselImProc.scala 113:21]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  stateReg = _RAND_0[1:0];
  _RAND_1 = {1{`RANDOM}};
  dataReg = _RAND_1[23:0];
  _RAND_2 = {1{`RANDOM}};
  shadowReg = _RAND_2[23:0];
  _RAND_3 = {1{`RANDOM}};
  userReg = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  shadowUserReg = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  lastReg = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  shadowLastReg = _RAND_6[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      stateReg <= 2'h0;
    end else if (_T) begin
      if (io_enq_valid) begin
        stateReg <= 2'h1;
      end
    end else if (_T_1) begin
      if (_T_3) begin
        stateReg <= 2'h0;
      end else if (_T_4) begin
        stateReg <= 2'h1;
      end else if (_T_6) begin
        stateReg <= 2'h2;
      end
    end else if (_T_7) begin
      if (io_deq_ready) begin
        stateReg <= 2'h1;
      end
    end else if (_T_8) begin
      stateReg <= 2'h0;
    end
    if (_T) begin
      if (io_enq_valid) begin
        dataReg <= io_enq_bits;
      end
    end else if (_T_1) begin
      if (!(_T_3)) begin
        if (_T_4) begin
          dataReg <= io_enq_bits;
        end
      end
    end else if (_T_7) begin
      if (io_deq_ready) begin
        dataReg <= shadowReg;
      end
    end
    if (!(_T)) begin
      if (_T_1) begin
        if (!(_T_3)) begin
          if (!(_T_4)) begin
            if (_T_6) begin
              shadowReg <= io_enq_bits;
            end
          end
        end
      end
    end
    if (_T) begin
      userReg <= io_enq_user;
    end else if (_T_1) begin
      if (_T_3) begin
        userReg <= io_enq_user;
      end else if (_T_4) begin
        userReg <= io_enq_user;
      end
    end else if (_T_7) begin
      if (io_deq_ready) begin
        userReg <= shadowUserReg;
      end
    end
    if (!(_T)) begin
      if (_T_1) begin
        if (!(_T_3)) begin
          if (!(_T_4)) begin
            if (_T_6) begin
              shadowUserReg <= io_enq_user;
            end
          end
        end
      end
    end
    if (_T) begin
      if (io_enq_valid) begin
        lastReg <= io_enq_last;
      end
    end else if (_T_1) begin
      if (!(_T_3)) begin
        if (_T_4) begin
          lastReg <= io_enq_last;
        end
      end
    end else if (_T_7) begin
      if (io_deq_ready) begin
        lastReg <= shadowLastReg;
      end
    end
    if (!(_T)) begin
      if (_T_1) begin
        if (!(_T_3)) begin
          if (!(_T_4)) begin
            if (_T_6) begin
              shadowLastReg <= io_enq_last;
            end
          end
        end
      end
    end
  end
endmodule
module ChiselImProc(
  input          clock,
  input          reset,
  output         io_enq_ready,
  input          io_enq_valid,
  input  [23:0]  io_enq_bits,
  input          io_enq_user,
  input          io_enq_last,
  input          io_deq_ready,
  output         io_deq_valid,
  output [23:0]  io_deq_bits,
  output         io_deq_user,
  output         io_deq_last,
  output [31:0]  io_dport,
  output [31:0]  io_dport2,
  output [15:0]  io_tdata,
  output [199:0] io_tdata2,
  output         io_tvalid,
  output         io_tready
);
  wire  RGB2GrayFilter_clock; // @[ChiselImProc.scala 503:16]
  wire  RGB2GrayFilter_reset; // @[ChiselImProc.scala 503:16]
  wire  RGB2GrayFilter_io_enq_ready; // @[ChiselImProc.scala 503:16]
  wire  RGB2GrayFilter_io_enq_valid; // @[ChiselImProc.scala 503:16]
  wire [23:0] RGB2GrayFilter_io_enq_bits; // @[ChiselImProc.scala 503:16]
  wire  RGB2GrayFilter_io_enq_user; // @[ChiselImProc.scala 503:16]
  wire  RGB2GrayFilter_io_enq_last; // @[ChiselImProc.scala 503:16]
  wire  RGB2GrayFilter_io_deq_ready; // @[ChiselImProc.scala 503:16]
  wire  RGB2GrayFilter_io_deq_valid; // @[ChiselImProc.scala 503:16]
  wire [23:0] RGB2GrayFilter_io_deq_bits; // @[ChiselImProc.scala 503:16]
  wire  RGB2GrayFilter_io_deq_user; // @[ChiselImProc.scala 503:16]
  wire  RGB2GrayFilter_io_deq_last; // @[ChiselImProc.scala 503:16]
  wire [8:0] RGB2GrayFilter_xcounter_0; // @[ChiselImProc.scala 503:16]
  wire [8:0] RGB2GrayFilter_ycounter_0; // @[ChiselImProc.scala 503:16]
  wire  GaussianBlurFilter_clock; // @[ChiselImProc.scala 505:16]
  wire  GaussianBlurFilter_reset; // @[ChiselImProc.scala 505:16]
  wire  GaussianBlurFilter_io__enq_ready; // @[ChiselImProc.scala 505:16]
  wire  GaussianBlurFilter_io__enq_valid; // @[ChiselImProc.scala 505:16]
  wire [7:0] GaussianBlurFilter_io__enq_bits; // @[ChiselImProc.scala 505:16]
  wire  GaussianBlurFilter_io__enq_user; // @[ChiselImProc.scala 505:16]
  wire  GaussianBlurFilter_io__enq_last; // @[ChiselImProc.scala 505:16]
  wire  GaussianBlurFilter_io__deq_ready; // @[ChiselImProc.scala 505:16]
  wire  GaussianBlurFilter_io__deq_valid; // @[ChiselImProc.scala 505:16]
  wire [7:0] GaussianBlurFilter_io__deq_bits; // @[ChiselImProc.scala 505:16]
  wire  GaussianBlurFilter_io__deq_user; // @[ChiselImProc.scala 505:16]
  wire  GaussianBlurFilter_io__deq_last; // @[ChiselImProc.scala 505:16]
  wire  GaussianBlurFilter_io_deq_ready; // @[ChiselImProc.scala 505:16]
  wire  GaussianBlurFilter_io_deq_valid; // @[ChiselImProc.scala 505:16]
  wire [71:0] GaussianBlurFilter__T_805_0; // @[ChiselImProc.scala 505:16]
  wire [15:0] GaussianBlurFilter_io_output; // @[ChiselImProc.scala 505:16]
  wire  SobelAndNonMaxSupressionFilter_clock; // @[ChiselImProc.scala 508:16]
  wire  SobelAndNonMaxSupressionFilter_reset; // @[ChiselImProc.scala 508:16]
  wire  SobelAndNonMaxSupressionFilter_io_enq_ready; // @[ChiselImProc.scala 508:16]
  wire  SobelAndNonMaxSupressionFilter_io_enq_valid; // @[ChiselImProc.scala 508:16]
  wire [7:0] SobelAndNonMaxSupressionFilter_io_enq_bits; // @[ChiselImProc.scala 508:16]
  wire  SobelAndNonMaxSupressionFilter_io_enq_user; // @[ChiselImProc.scala 508:16]
  wire  SobelAndNonMaxSupressionFilter_io_enq_last; // @[ChiselImProc.scala 508:16]
  wire  SobelAndNonMaxSupressionFilter_io_deq_ready; // @[ChiselImProc.scala 508:16]
  wire  SobelAndNonMaxSupressionFilter_io_deq_valid; // @[ChiselImProc.scala 508:16]
  wire [7:0] SobelAndNonMaxSupressionFilter_io_deq_bits; // @[ChiselImProc.scala 508:16]
  wire  SobelAndNonMaxSupressionFilter_io_deq_user; // @[ChiselImProc.scala 508:16]
  wire  SobelAndNonMaxSupressionFilter_io_deq_last; // @[ChiselImProc.scala 508:16]
  wire  ZeroPadding_clock; // @[ChiselImProc.scala 512:16]
  wire  ZeroPadding_reset; // @[ChiselImProc.scala 512:16]
  wire  ZeroPadding_io_enq_ready; // @[ChiselImProc.scala 512:16]
  wire  ZeroPadding_io_enq_valid; // @[ChiselImProc.scala 512:16]
  wire [7:0] ZeroPadding_io_enq_bits; // @[ChiselImProc.scala 512:16]
  wire  ZeroPadding_io_enq_user; // @[ChiselImProc.scala 512:16]
  wire  ZeroPadding_io_enq_last; // @[ChiselImProc.scala 512:16]
  wire  ZeroPadding_io_deq_ready; // @[ChiselImProc.scala 512:16]
  wire  ZeroPadding_io_deq_valid; // @[ChiselImProc.scala 512:16]
  wire [7:0] ZeroPadding_io_deq_bits; // @[ChiselImProc.scala 512:16]
  wire  ZeroPadding_io_deq_user; // @[ChiselImProc.scala 512:16]
  wire  ZeroPadding_io_deq_last; // @[ChiselImProc.scala 512:16]
  wire  HystThreshold_clock; // @[ChiselImProc.scala 515:16]
  wire  HystThreshold_reset; // @[ChiselImProc.scala 515:16]
  wire  HystThreshold_io_enq_ready; // @[ChiselImProc.scala 515:16]
  wire  HystThreshold_io_enq_valid; // @[ChiselImProc.scala 515:16]
  wire [7:0] HystThreshold_io_enq_bits; // @[ChiselImProc.scala 515:16]
  wire  HystThreshold_io_enq_user; // @[ChiselImProc.scala 515:16]
  wire  HystThreshold_io_enq_last; // @[ChiselImProc.scala 515:16]
  wire  HystThreshold_io_deq_ready; // @[ChiselImProc.scala 515:16]
  wire  HystThreshold_io_deq_valid; // @[ChiselImProc.scala 515:16]
  wire [7:0] HystThreshold_io_deq_bits; // @[ChiselImProc.scala 515:16]
  wire  HystThreshold_io_deq_user; // @[ChiselImProc.scala 515:16]
  wire  HystThreshold_io_deq_last; // @[ChiselImProc.scala 515:16]
  wire  HystThresholdComp_clock; // @[ChiselImProc.scala 518:16]
  wire  HystThresholdComp_reset; // @[ChiselImProc.scala 518:16]
  wire  HystThresholdComp_io_enq_ready; // @[ChiselImProc.scala 518:16]
  wire  HystThresholdComp_io_enq_valid; // @[ChiselImProc.scala 518:16]
  wire [7:0] HystThresholdComp_io_enq_bits; // @[ChiselImProc.scala 518:16]
  wire  HystThresholdComp_io_enq_user; // @[ChiselImProc.scala 518:16]
  wire  HystThresholdComp_io_enq_last; // @[ChiselImProc.scala 518:16]
  wire  HystThresholdComp_io_deq_ready; // @[ChiselImProc.scala 518:16]
  wire  HystThresholdComp_io_deq_valid; // @[ChiselImProc.scala 518:16]
  wire [7:0] HystThresholdComp_io_deq_bits; // @[ChiselImProc.scala 518:16]
  wire  HystThresholdComp_io_deq_user; // @[ChiselImProc.scala 518:16]
  wire  HystThresholdComp_io_deq_last; // @[ChiselImProc.scala 518:16]
  wire  Gray2RGBFilter_clock; // @[ChiselImProc.scala 521:16]
  wire  Gray2RGBFilter_reset; // @[ChiselImProc.scala 521:16]
  wire  Gray2RGBFilter_io_enq_ready; // @[ChiselImProc.scala 521:16]
  wire  Gray2RGBFilter_io_enq_valid; // @[ChiselImProc.scala 521:16]
  wire [23:0] Gray2RGBFilter_io_enq_bits; // @[ChiselImProc.scala 521:16]
  wire  Gray2RGBFilter_io_enq_user; // @[ChiselImProc.scala 521:16]
  wire  Gray2RGBFilter_io_enq_last; // @[ChiselImProc.scala 521:16]
  wire  Gray2RGBFilter_io_deq_ready; // @[ChiselImProc.scala 521:16]
  wire  Gray2RGBFilter_io_deq_valid; // @[ChiselImProc.scala 521:16]
  wire [23:0] Gray2RGBFilter_io_deq_bits; // @[ChiselImProc.scala 521:16]
  wire  Gray2RGBFilter_io_deq_user; // @[ChiselImProc.scala 521:16]
  wire  Gray2RGBFilter_io_deq_last; // @[ChiselImProc.scala 521:16]
  wire [71:0] tdata2_0 = GaussianBlurFilter__T_805_0;
  wire [8:0] uniqueId2 = RGB2GrayFilter_ycounter_0;
  wire [8:0] uniqueId = RGB2GrayFilter_xcounter_0;
  RGB2GrayFilter RGB2GrayFilter ( // @[ChiselImProc.scala 503:16]
    .clock(RGB2GrayFilter_clock),
    .reset(RGB2GrayFilter_reset),
    .io_enq_ready(RGB2GrayFilter_io_enq_ready),
    .io_enq_valid(RGB2GrayFilter_io_enq_valid),
    .io_enq_bits(RGB2GrayFilter_io_enq_bits),
    .io_enq_user(RGB2GrayFilter_io_enq_user),
    .io_enq_last(RGB2GrayFilter_io_enq_last),
    .io_deq_ready(RGB2GrayFilter_io_deq_ready),
    .io_deq_valid(RGB2GrayFilter_io_deq_valid),
    .io_deq_bits(RGB2GrayFilter_io_deq_bits),
    .io_deq_user(RGB2GrayFilter_io_deq_user),
    .io_deq_last(RGB2GrayFilter_io_deq_last),
    .xcounter_0(RGB2GrayFilter_xcounter_0),
    .ycounter_0(RGB2GrayFilter_ycounter_0)
  );
  GaussianBlurFilter GaussianBlurFilter ( // @[ChiselImProc.scala 505:16]
    .clock(GaussianBlurFilter_clock),
    .reset(GaussianBlurFilter_reset),
    .io__enq_ready(GaussianBlurFilter_io__enq_ready),
    .io__enq_valid(GaussianBlurFilter_io__enq_valid),
    .io__enq_bits(GaussianBlurFilter_io__enq_bits),
    .io__enq_user(GaussianBlurFilter_io__enq_user),
    .io__enq_last(GaussianBlurFilter_io__enq_last),
    .io__deq_ready(GaussianBlurFilter_io__deq_ready),
    .io__deq_valid(GaussianBlurFilter_io__deq_valid),
    .io__deq_bits(GaussianBlurFilter_io__deq_bits),
    .io__deq_user(GaussianBlurFilter_io__deq_user),
    .io__deq_last(GaussianBlurFilter_io__deq_last),
    .io_deq_ready(GaussianBlurFilter_io_deq_ready),
    .io_deq_valid(GaussianBlurFilter_io_deq_valid),
    ._T_805_0(GaussianBlurFilter__T_805_0),
    .io_output(GaussianBlurFilter_io_output)
  );
  SobelAndNonMaxSupressionFilter SobelAndNonMaxSupressionFilter ( // @[ChiselImProc.scala 508:16]
    .clock(SobelAndNonMaxSupressionFilter_clock),
    .reset(SobelAndNonMaxSupressionFilter_reset),
    .io_enq_ready(SobelAndNonMaxSupressionFilter_io_enq_ready),
    .io_enq_valid(SobelAndNonMaxSupressionFilter_io_enq_valid),
    .io_enq_bits(SobelAndNonMaxSupressionFilter_io_enq_bits),
    .io_enq_user(SobelAndNonMaxSupressionFilter_io_enq_user),
    .io_enq_last(SobelAndNonMaxSupressionFilter_io_enq_last),
    .io_deq_ready(SobelAndNonMaxSupressionFilter_io_deq_ready),
    .io_deq_valid(SobelAndNonMaxSupressionFilter_io_deq_valid),
    .io_deq_bits(SobelAndNonMaxSupressionFilter_io_deq_bits),
    .io_deq_user(SobelAndNonMaxSupressionFilter_io_deq_user),
    .io_deq_last(SobelAndNonMaxSupressionFilter_io_deq_last)
  );
  ZeroPadding ZeroPadding ( // @[ChiselImProc.scala 512:16]
    .clock(ZeroPadding_clock),
    .reset(ZeroPadding_reset),
    .io_enq_ready(ZeroPadding_io_enq_ready),
    .io_enq_valid(ZeroPadding_io_enq_valid),
    .io_enq_bits(ZeroPadding_io_enq_bits),
    .io_enq_user(ZeroPadding_io_enq_user),
    .io_enq_last(ZeroPadding_io_enq_last),
    .io_deq_ready(ZeroPadding_io_deq_ready),
    .io_deq_valid(ZeroPadding_io_deq_valid),
    .io_deq_bits(ZeroPadding_io_deq_bits),
    .io_deq_user(ZeroPadding_io_deq_user),
    .io_deq_last(ZeroPadding_io_deq_last)
  );
  HystThreshold HystThreshold ( // @[ChiselImProc.scala 515:16]
    .clock(HystThreshold_clock),
    .reset(HystThreshold_reset),
    .io_enq_ready(HystThreshold_io_enq_ready),
    .io_enq_valid(HystThreshold_io_enq_valid),
    .io_enq_bits(HystThreshold_io_enq_bits),
    .io_enq_user(HystThreshold_io_enq_user),
    .io_enq_last(HystThreshold_io_enq_last),
    .io_deq_ready(HystThreshold_io_deq_ready),
    .io_deq_valid(HystThreshold_io_deq_valid),
    .io_deq_bits(HystThreshold_io_deq_bits),
    .io_deq_user(HystThreshold_io_deq_user),
    .io_deq_last(HystThreshold_io_deq_last)
  );
  HystThresholdComp HystThresholdComp ( // @[ChiselImProc.scala 518:16]
    .clock(HystThresholdComp_clock),
    .reset(HystThresholdComp_reset),
    .io_enq_ready(HystThresholdComp_io_enq_ready),
    .io_enq_valid(HystThresholdComp_io_enq_valid),
    .io_enq_bits(HystThresholdComp_io_enq_bits),
    .io_enq_user(HystThresholdComp_io_enq_user),
    .io_enq_last(HystThresholdComp_io_enq_last),
    .io_deq_ready(HystThresholdComp_io_deq_ready),
    .io_deq_valid(HystThresholdComp_io_deq_valid),
    .io_deq_bits(HystThresholdComp_io_deq_bits),
    .io_deq_user(HystThresholdComp_io_deq_user),
    .io_deq_last(HystThresholdComp_io_deq_last)
  );
  Gray2RGBFilter Gray2RGBFilter ( // @[ChiselImProc.scala 521:16]
    .clock(Gray2RGBFilter_clock),
    .reset(Gray2RGBFilter_reset),
    .io_enq_ready(Gray2RGBFilter_io_enq_ready),
    .io_enq_valid(Gray2RGBFilter_io_enq_valid),
    .io_enq_bits(Gray2RGBFilter_io_enq_bits),
    .io_enq_user(Gray2RGBFilter_io_enq_user),
    .io_enq_last(Gray2RGBFilter_io_enq_last),
    .io_deq_ready(Gray2RGBFilter_io_deq_ready),
    .io_deq_valid(Gray2RGBFilter_io_deq_valid),
    .io_deq_bits(Gray2RGBFilter_io_deq_bits),
    .io_deq_user(Gray2RGBFilter_io_deq_user),
    .io_deq_last(Gray2RGBFilter_io_deq_last)
  );
  assign io_enq_ready = RGB2GrayFilter_io_enq_ready; // @[ChiselImProc.scala 532:12]
  assign io_deq_valid = Gray2RGBFilter_io_deq_valid; // @[ChiselImProc.scala 534:12]
  assign io_deq_bits = Gray2RGBFilter_io_deq_bits; // @[ChiselImProc.scala 534:12]
  assign io_deq_user = Gray2RGBFilter_io_deq_user; // @[ChiselImProc.scala 534:12]
  assign io_deq_last = Gray2RGBFilter_io_deq_last; // @[ChiselImProc.scala 534:12]
  assign io_dport = {{23'd0}, uniqueId}; // @[ChiselImProc.scala 560:14]
  assign io_dport2 = {{23'd0}, uniqueId2}; // @[ChiselImProc.scala 561:15]
  assign io_tdata = GaussianBlurFilter_io_output; // @[ChiselImProc.scala 562:14]
  assign io_tdata2 = {{128'd0}, tdata2_0}; // @[ChiselImProc.scala 565:15]
  assign io_tvalid = GaussianBlurFilter_io_deq_valid; // @[ChiselImProc.scala 563:15]
  assign io_tready = GaussianBlurFilter_io_deq_ready; // @[ChiselImProc.scala 564:15]
  assign RGB2GrayFilter_clock = clock;
  assign RGB2GrayFilter_reset = reset;
  assign RGB2GrayFilter_io_enq_valid = io_enq_valid; // @[ChiselImProc.scala 532:12]
  assign RGB2GrayFilter_io_enq_bits = io_enq_bits; // @[ChiselImProc.scala 532:12]
  assign RGB2GrayFilter_io_enq_user = io_enq_user; // @[ChiselImProc.scala 532:12]
  assign RGB2GrayFilter_io_enq_last = io_enq_last; // @[ChiselImProc.scala 532:12]
  assign RGB2GrayFilter_io_deq_ready = GaussianBlurFilter_io__enq_ready; // @[ChiselImProc.scala 529:30]
  assign GaussianBlurFilter_clock = clock;
  assign GaussianBlurFilter_reset = reset;
  assign GaussianBlurFilter_io__enq_valid = RGB2GrayFilter_io_deq_valid; // @[ChiselImProc.scala 529:30]
  assign GaussianBlurFilter_io__enq_bits = RGB2GrayFilter_io_deq_bits[7:0]; // @[ChiselImProc.scala 529:30]
  assign GaussianBlurFilter_io__enq_user = RGB2GrayFilter_io_deq_user; // @[ChiselImProc.scala 529:30]
  assign GaussianBlurFilter_io__enq_last = RGB2GrayFilter_io_deq_last; // @[ChiselImProc.scala 529:30]
  assign GaussianBlurFilter_io__deq_ready = SobelAndNonMaxSupressionFilter_io_enq_ready; // @[ChiselImProc.scala 529:30]
  assign SobelAndNonMaxSupressionFilter_clock = clock;
  assign SobelAndNonMaxSupressionFilter_reset = reset;
  assign SobelAndNonMaxSupressionFilter_io_enq_valid = GaussianBlurFilter_io__deq_valid; // @[ChiselImProc.scala 529:30]
  assign SobelAndNonMaxSupressionFilter_io_enq_bits = GaussianBlurFilter_io__deq_bits; // @[ChiselImProc.scala 529:30]
  assign SobelAndNonMaxSupressionFilter_io_enq_user = GaussianBlurFilter_io__deq_user; // @[ChiselImProc.scala 529:30]
  assign SobelAndNonMaxSupressionFilter_io_enq_last = GaussianBlurFilter_io__deq_last; // @[ChiselImProc.scala 529:30]
  assign SobelAndNonMaxSupressionFilter_io_deq_ready = ZeroPadding_io_enq_ready; // @[ChiselImProc.scala 529:30]
  assign ZeroPadding_clock = clock;
  assign ZeroPadding_reset = reset;
  assign ZeroPadding_io_enq_valid = SobelAndNonMaxSupressionFilter_io_deq_valid; // @[ChiselImProc.scala 529:30]
  assign ZeroPadding_io_enq_bits = SobelAndNonMaxSupressionFilter_io_deq_bits; // @[ChiselImProc.scala 529:30]
  assign ZeroPadding_io_enq_user = SobelAndNonMaxSupressionFilter_io_deq_user; // @[ChiselImProc.scala 529:30]
  assign ZeroPadding_io_enq_last = SobelAndNonMaxSupressionFilter_io_deq_last; // @[ChiselImProc.scala 529:30]
  assign ZeroPadding_io_deq_ready = HystThreshold_io_enq_ready; // @[ChiselImProc.scala 529:30]
  assign HystThreshold_clock = clock;
  assign HystThreshold_reset = reset;
  assign HystThreshold_io_enq_valid = ZeroPadding_io_deq_valid; // @[ChiselImProc.scala 529:30]
  assign HystThreshold_io_enq_bits = ZeroPadding_io_deq_bits; // @[ChiselImProc.scala 529:30]
  assign HystThreshold_io_enq_user = ZeroPadding_io_deq_user; // @[ChiselImProc.scala 529:30]
  assign HystThreshold_io_enq_last = ZeroPadding_io_deq_last; // @[ChiselImProc.scala 529:30]
  assign HystThreshold_io_deq_ready = HystThresholdComp_io_enq_ready; // @[ChiselImProc.scala 529:30]
  assign HystThresholdComp_clock = clock;
  assign HystThresholdComp_reset = reset;
  assign HystThresholdComp_io_enq_valid = HystThreshold_io_deq_valid; // @[ChiselImProc.scala 529:30]
  assign HystThresholdComp_io_enq_bits = HystThreshold_io_deq_bits; // @[ChiselImProc.scala 529:30]
  assign HystThresholdComp_io_enq_user = HystThreshold_io_deq_user; // @[ChiselImProc.scala 529:30]
  assign HystThresholdComp_io_enq_last = HystThreshold_io_deq_last; // @[ChiselImProc.scala 529:30]
  assign HystThresholdComp_io_deq_ready = Gray2RGBFilter_io_enq_ready; // @[ChiselImProc.scala 529:30]
  assign Gray2RGBFilter_clock = clock;
  assign Gray2RGBFilter_reset = reset;
  assign Gray2RGBFilter_io_enq_valid = HystThresholdComp_io_deq_valid; // @[ChiselImProc.scala 529:30]
  assign Gray2RGBFilter_io_enq_bits = {{16'd0}, HystThresholdComp_io_deq_bits}; // @[ChiselImProc.scala 529:30]
  assign Gray2RGBFilter_io_enq_user = HystThresholdComp_io_deq_user; // @[ChiselImProc.scala 529:30]
  assign Gray2RGBFilter_io_enq_last = HystThresholdComp_io_deq_last; // @[ChiselImProc.scala 529:30]
  assign Gray2RGBFilter_io_deq_ready = io_deq_ready; // @[ChiselImProc.scala 534:12]
endmodule

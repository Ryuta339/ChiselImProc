module SqrtExtractionUInt(
  input         clock,
  input         reset,
  input  [15:0] io_z,
  output [7:0]  io_q
);
  wire [16:0] zj_7 = {1'h0,io_z[15:14],14'h0}; // @[Cat.scala 29:58]
  wire [2:0] _T_5 = zj_7[16:14] - 3'h1; // @[Sqrt.scala 54:77]
  wire [16:0] rj_7 = {_T_5,14'h0}; // @[Cat.scala 29:58]
  wire  qSub_7 = ~rj_7[16]; // @[Sqrt.scala 55:27]
  wire [13:0] _T_14 = {io_z[13:12],12'h0}; // @[Cat.scala 29:58]
  wire [16:0] zj_6 = {{3'd0}, _T_14}; // @[Sqrt.scala 47:19 Sqrt.scala 59:19 Sqrt.scala 61:19 Sqrt.scala 64:19]
  wire [2:0] _T_18 = {qSub_7,2'h1}; // @[Cat.scala 29:58]
  wire [4:0] _GEN_7 = {{2'd0}, _T_18}; // @[Sqrt.scala 66:54]
  wire [4:0] _T_20 = zj_6[16:12] - _GEN_7; // @[Sqrt.scala 66:54]
  wire [16:0] rj_6 = {_T_20,12'h0}; // @[Cat.scala 29:58]
  wire  qSub_6 = ~rj_6[16]; // @[Sqrt.scala 72:20]
  wire [11:0] _T_29 = {io_z[11:10],10'h0}; // @[Cat.scala 29:58]
  wire [16:0] zj_5 = {{5'd0}, _T_29}; // @[Sqrt.scala 47:19 Sqrt.scala 59:19 Sqrt.scala 61:19 Sqrt.scala 64:19]
  wire [3:0] _T_34 = {qSub_7,qSub_6,2'h1}; // @[Cat.scala 29:58]
  wire [5:0] _GEN_8 = {{2'd0}, _T_34}; // @[Sqrt.scala 66:54]
  wire [5:0] _T_36 = zj_5[15:10] - _GEN_8; // @[Sqrt.scala 66:54]
  wire [15:0] _T_37 = {_T_36,10'h0}; // @[Cat.scala 29:58]
  wire [16:0] rj_5 = {{1'd0}, _T_37}; // @[Sqrt.scala 48:19 Sqrt.scala 66:19]
  wire  qSub_5 = ~rj_5[15]; // @[Sqrt.scala 72:20]
  wire [9:0] _T_45 = {io_z[9:8],8'h0}; // @[Cat.scala 29:58]
  wire [16:0] zj_4 = {{7'd0}, _T_45}; // @[Sqrt.scala 47:19 Sqrt.scala 59:19 Sqrt.scala 61:19 Sqrt.scala 64:19]
  wire [4:0] _T_51 = {qSub_7,qSub_6,qSub_5,2'h1}; // @[Cat.scala 29:58]
  wire [6:0] _GEN_9 = {{2'd0}, _T_51}; // @[Sqrt.scala 66:54]
  wire [6:0] _T_53 = zj_4[14:8] - _GEN_9; // @[Sqrt.scala 66:54]
  wire [14:0] _T_54 = {_T_53,8'h0}; // @[Cat.scala 29:58]
  wire [16:0] rj_4 = {{2'd0}, _T_54}; // @[Sqrt.scala 48:19 Sqrt.scala 66:19]
  wire  qSub_4 = ~rj_4[14]; // @[Sqrt.scala 72:20]
  wire [7:0] _T_62 = {io_z[7:6],6'h0}; // @[Cat.scala 29:58]
  wire [16:0] zj_3 = {{9'd0}, _T_62}; // @[Sqrt.scala 47:19 Sqrt.scala 59:19 Sqrt.scala 61:19 Sqrt.scala 64:19]
  wire [3:0] _T_68 = {qSub_7,qSub_6,qSub_5,qSub_4}; // @[Sqrt.scala 66:67]
  wire [5:0] _T_69 = {qSub_7,qSub_6,qSub_5,qSub_4,2'h1}; // @[Cat.scala 29:58]
  wire [7:0] _GEN_10 = {{2'd0}, _T_69}; // @[Sqrt.scala 66:54]
  wire [7:0] _T_71 = zj_3[13:6] - _GEN_10; // @[Sqrt.scala 66:54]
  wire [13:0] _T_72 = {_T_71,6'h0}; // @[Cat.scala 29:58]
  wire [16:0] rj_3 = {{3'd0}, _T_72}; // @[Sqrt.scala 48:19 Sqrt.scala 66:19]
  wire  qSub_3 = ~rj_3[13]; // @[Sqrt.scala 72:20]
  wire [5:0] _T_80 = {io_z[5:4],4'h0}; // @[Cat.scala 29:58]
  wire [16:0] zj_2 = {{11'd0}, _T_80}; // @[Sqrt.scala 47:19 Sqrt.scala 59:19 Sqrt.scala 61:19 Sqrt.scala 64:19]
  wire [6:0] _T_88 = {qSub_7,qSub_6,qSub_5,qSub_4,qSub_3,2'h1}; // @[Cat.scala 29:58]
  wire [8:0] _GEN_11 = {{2'd0}, _T_88}; // @[Sqrt.scala 66:54]
  wire [8:0] _T_90 = zj_2[12:4] - _GEN_11; // @[Sqrt.scala 66:54]
  wire [12:0] _T_91 = {_T_90,4'h0}; // @[Cat.scala 29:58]
  wire [16:0] rj_2 = {{4'd0}, _T_91}; // @[Sqrt.scala 48:19 Sqrt.scala 66:19]
  wire  qSub_2 = ~rj_2[12]; // @[Sqrt.scala 72:20]
  wire [3:0] _T_99 = {io_z[3:2],2'h0}; // @[Cat.scala 29:58]
  wire [16:0] zj_1 = {{13'd0}, _T_99}; // @[Sqrt.scala 47:19 Sqrt.scala 59:19 Sqrt.scala 61:19 Sqrt.scala 64:19]
  wire [7:0] _T_108 = {qSub_7,qSub_6,qSub_5,qSub_4,qSub_3,qSub_2,2'h1}; // @[Cat.scala 29:58]
  wire [9:0] _GEN_12 = {{2'd0}, _T_108}; // @[Sqrt.scala 66:54]
  wire [9:0] _T_110 = zj_1[11:2] - _GEN_12; // @[Sqrt.scala 66:54]
  wire [11:0] _T_111 = {_T_110,2'h0}; // @[Cat.scala 29:58]
  wire [16:0] rj_1 = {{5'd0}, _T_111}; // @[Sqrt.scala 48:19 Sqrt.scala 66:19]
  wire  qSub_1 = ~rj_1[11]; // @[Sqrt.scala 72:20]
  wire [16:0] zj_0 = {{15'd0}, io_z[1:0]}; // @[Sqrt.scala 47:19 Sqrt.scala 59:19 Sqrt.scala 61:19 Sqrt.scala 68:19]
  wire [8:0] _T_128 = {qSub_7,qSub_6,qSub_5,qSub_4,qSub_3,qSub_2,qSub_1,2'h1}; // @[Cat.scala 29:58]
  wire [10:0] _GEN_13 = {{2'd0}, _T_128}; // @[Sqrt.scala 70:49]
  wire [10:0] _T_130 = zj_0[10:0] - _GEN_13; // @[Sqrt.scala 70:49]
  wire [16:0] rj_0 = {{6'd0}, _T_130}; // @[Sqrt.scala 48:19 Sqrt.scala 70:19]
  wire  qSub_0 = ~rj_0[10]; // @[Sqrt.scala 72:20]
  wire [3:0] _T_135 = {qSub_3,qSub_2,qSub_1,qSub_0}; // @[Sqrt.scala 75:18]
  assign io_q = {_T_68,_T_135}; // @[Sqrt.scala 75:10]
endmodule

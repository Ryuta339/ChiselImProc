// axi4.ImProcMain1913971855
// 2020/12/02 13:00

module RGB2GrayFilter(
  input         clock,
  input         reset,
  output        io_enq_ready,
  input         io_enq_valid,
  input  [23:0] io_enq_bits,
  input         io_enq_user,
  input         io_enq_last,
  input         io_deq_ready,
  output        io_deq_valid,
  output [23:0] io_deq_bits,
  output        io_deq_user,
  output        io_deq_last
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
`endif // RANDOMIZE_REG_INIT
  reg [1:0] stateReg; // @[ChiselImProc.scala 56:28]
  reg [23:0] dataReg; // @[ChiselImProc.scala 58:23]
  reg [23:0] shadowReg; // @[ChiselImProc.scala 60:25]
  reg  userReg; // @[ChiselImProc.scala 61:23]
  reg  shadowUserReg; // @[ChiselImProc.scala 62:29]
  reg  lastReg; // @[ChiselImProc.scala 63:23]
  reg  shadowLastReg; // @[ChiselImProc.scala 64:29]
  wire  _T = 2'h0 == stateReg; // @[Conditional.scala 37:30]
  wire  _T_1 = 2'h1 == stateReg; // @[Conditional.scala 37:30]
  wire  _T_2 = ~io_enq_valid; // @[ChiselImProc.scala 78:39]
  wire  _T_3 = io_deq_ready & _T_2; // @[ChiselImProc.scala 78:36]
  wire  _T_4 = io_deq_ready & io_enq_valid; // @[ChiselImProc.scala 81:42]
  wire  _T_5 = ~io_deq_ready; // @[ChiselImProc.scala 86:29]
  wire  _T_6 = _T_5 & io_enq_valid; // @[ChiselImProc.scala 86:43]
  wire  _T_7 = 2'h2 == stateReg; // @[Conditional.scala 37:30]
  wire  _T_8 = 2'h3 == stateReg; // @[Conditional.scala 37:30]
  wire  _T_9 = stateReg == 2'h0; // @[ChiselImProc.scala 110:35]
  wire  _T_10 = stateReg == 2'h1; // @[ChiselImProc.scala 110:57]
  wire  _T_11 = _T_9 | _T_10; // @[ChiselImProc.scala 110:45]
  wire  _T_12 = stateReg == 2'h3; // @[ChiselImProc.scala 110:77]
  wire  _T_15 = stateReg == 2'h2; // @[ChiselImProc.scala 111:55]
  wire [23:0] _T_17 = dataReg & 24'hff; // @[ChiselImProc.scala 163:36]
  wire [37:0] _T_18 = 24'h24dd * _T_17; // @[ChiselImProc.scala 163:25]
  wire [23:0] _T_19 = dataReg & 24'hff00; // @[ChiselImProc.scala 164:33]
  wire [23:0] _T_20 = {{8'd0}, _T_19[23:8]}; // @[ChiselImProc.scala 164:47]
  wire [39:0] _T_21 = 24'h9645 * _T_20; // @[ChiselImProc.scala 164:21]
  wire [39:0] _GEN_45 = {{2'd0}, _T_18}; // @[ChiselImProc.scala 163:50]
  wire [39:0] _T_23 = _GEN_45 + _T_21; // @[ChiselImProc.scala 163:50]
  wire [23:0] _T_24 = dataReg & 24'hff0000; // @[ChiselImProc.scala 165:33]
  wire [23:0] _T_25 = {{16'd0}, _T_24[23:16]}; // @[ChiselImProc.scala 165:47]
  wire [38:0] _T_26 = 24'h4c8b * _T_25; // @[ChiselImProc.scala 165:21]
  wire [39:0] _GEN_47 = {{1'd0}, _T_26}; // @[ChiselImProc.scala 164:55]
  wire [39:0] _T_28 = _T_23 + _GEN_47; // @[ChiselImProc.scala 164:55]
  wire [31:0] pixGray = _T_28[31:0]; // @[ChiselImProc.scala 160:24 ChiselImProc.scala 163:13]
  wire [31:0] _T_29 = {{16'd0}, pixGray[31:16]}; // @[ChiselImProc.scala 167:24]
  wire [15:0] rolled = _T_29[15:0]; // @[ChiselImProc.scala 161:23 ChiselImProc.scala 167:12]
  wire  _T_30 = rolled > 16'hff; // @[ChiselImProc.scala 168:32]
  wire [15:0] _T_31 = _T_30 ? 16'hff : rolled; // @[ChiselImProc.scala 168:24]
  assign io_enq_ready = _T_11 | _T_12; // @[ChiselImProc.scala 110:22]
  assign io_deq_valid = _T_10 | _T_15; // @[ChiselImProc.scala 111:22]
  assign io_deq_bits = {{8'd0}, _T_31}; // @[ChiselImProc.scala 168:17]
  assign io_deq_user = userReg; // @[ChiselImProc.scala 138:17 ChiselImProc.scala 108:21]
  assign io_deq_last = lastReg; // @[ChiselImProc.scala 137:17 ChiselImProc.scala 107:21]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  stateReg = _RAND_0[1:0];
  _RAND_1 = {1{`RANDOM}};
  dataReg = _RAND_1[23:0];
  _RAND_2 = {1{`RANDOM}};
  shadowReg = _RAND_2[23:0];
  _RAND_3 = {1{`RANDOM}};
  userReg = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  shadowUserReg = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  lastReg = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  shadowLastReg = _RAND_6[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      stateReg <= 2'h0;
    end else if (_T) begin
      if (io_enq_valid) begin
        stateReg <= 2'h1;
      end
    end else if (_T_1) begin
      if (_T_3) begin
        stateReg <= 2'h0;
      end else if (_T_4) begin
        stateReg <= 2'h1;
      end else if (_T_6) begin
        stateReg <= 2'h2;
      end
    end else if (_T_7) begin
      if (io_deq_ready) begin
        stateReg <= 2'h1;
      end
    end else if (_T_8) begin
      stateReg <= 2'h0;
    end
    if (_T) begin
      if (io_enq_valid) begin
        dataReg <= io_enq_bits;
      end
    end else if (_T_1) begin
      if (!(_T_3)) begin
        if (_T_4) begin
          dataReg <= io_enq_bits;
        end
      end
    end else if (_T_7) begin
      if (io_deq_ready) begin
        dataReg <= shadowReg;
      end
    end
    if (!(_T)) begin
      if (_T_1) begin
        if (!(_T_3)) begin
          if (!(_T_4)) begin
            if (_T_6) begin
              shadowReg <= io_enq_bits;
            end
          end
        end
      end
    end
    if (_T) begin
      userReg <= io_enq_user;
    end else if (_T_1) begin
      if (_T_3) begin
        userReg <= io_enq_user;
      end else if (_T_4) begin
        userReg <= io_enq_user;
      end
    end else if (_T_7) begin
      if (io_deq_ready) begin
        userReg <= shadowUserReg;
      end
    end
    if (!(_T)) begin
      if (_T_1) begin
        if (!(_T_3)) begin
          if (!(_T_4)) begin
            if (_T_6) begin
              shadowUserReg <= io_enq_user;
            end
          end
        end
      end
    end
    if (_T) begin
      if (io_enq_valid) begin
        lastReg <= io_enq_last;
      end
    end else if (_T_1) begin
      if (!(_T_3)) begin
        if (_T_4) begin
          lastReg <= io_enq_last;
        end
      end
    end else if (_T_7) begin
      if (io_deq_ready) begin
        lastReg <= shadowLastReg;
      end
    end
    if (!(_T)) begin
      if (_T_1) begin
        if (!(_T_3)) begin
          if (!(_T_4)) begin
            if (_T_6) begin
              shadowLastReg <= io_enq_last;
            end
          end
        end
      end
    end
  end
endmodule
module MulAdd(
  input  [7:0]  io_b_0,
  input  [7:0]  io_b_1,
  input  [7:0]  io_b_2,
  input  [7:0]  io_b_3,
  input  [7:0]  io_b_4,
  input  [7:0]  io_b_5,
  input  [7:0]  io_b_6,
  input  [7:0]  io_b_7,
  input  [7:0]  io_b_8,
  input  [7:0]  io_b_9,
  input  [7:0]  io_b_10,
  input  [7:0]  io_b_11,
  input  [7:0]  io_b_12,
  input  [7:0]  io_b_13,
  input  [7:0]  io_b_14,
  input  [7:0]  io_b_15,
  input  [7:0]  io_b_16,
  input  [7:0]  io_b_17,
  input  [7:0]  io_b_18,
  input  [7:0]  io_b_19,
  input  [7:0]  io_b_20,
  input  [7:0]  io_b_21,
  input  [7:0]  io_b_22,
  input  [7:0]  io_b_23,
  input  [7:0]  io_b_24,
  output [15:0] io_output
);
  wire [15:0] _T = 8'h1 * io_b_0; // @[ChiselImProc.scala 28:24]
  wire [16:0] _T_1 = {{1'd0}, _T}; // @[ChiselImProc.scala 28:13]
  wire [15:0] _T_3 = 8'h4 * io_b_1; // @[ChiselImProc.scala 28:24]
  wire [15:0] _T_5 = _T_1[15:0] + _T_3; // @[ChiselImProc.scala 28:13]
  wire [15:0] _T_6 = 8'h6 * io_b_2; // @[ChiselImProc.scala 28:24]
  wire [15:0] _T_8 = _T_5 + _T_6; // @[ChiselImProc.scala 28:13]
  wire [15:0] _T_9 = 8'h4 * io_b_3; // @[ChiselImProc.scala 28:24]
  wire [15:0] _T_11 = _T_8 + _T_9; // @[ChiselImProc.scala 28:13]
  wire [15:0] _T_12 = 8'h1 * io_b_4; // @[ChiselImProc.scala 28:24]
  wire [15:0] _T_14 = _T_11 + _T_12; // @[ChiselImProc.scala 28:13]
  wire [15:0] _T_15 = 8'h4 * io_b_5; // @[ChiselImProc.scala 28:24]
  wire [15:0] _T_17 = _T_14 + _T_15; // @[ChiselImProc.scala 28:13]
  wire [15:0] _T_18 = 8'h10 * io_b_6; // @[ChiselImProc.scala 28:24]
  wire [15:0] _T_20 = _T_17 + _T_18; // @[ChiselImProc.scala 28:13]
  wire [15:0] _T_21 = 8'h18 * io_b_7; // @[ChiselImProc.scala 28:24]
  wire [15:0] _T_23 = _T_20 + _T_21; // @[ChiselImProc.scala 28:13]
  wire [15:0] _T_24 = 8'h10 * io_b_8; // @[ChiselImProc.scala 28:24]
  wire [15:0] _T_26 = _T_23 + _T_24; // @[ChiselImProc.scala 28:13]
  wire [15:0] _T_27 = 8'h4 * io_b_9; // @[ChiselImProc.scala 28:24]
  wire [15:0] _T_29 = _T_26 + _T_27; // @[ChiselImProc.scala 28:13]
  wire [15:0] _T_30 = 8'h6 * io_b_10; // @[ChiselImProc.scala 28:24]
  wire [15:0] _T_32 = _T_29 + _T_30; // @[ChiselImProc.scala 28:13]
  wire [15:0] _T_33 = 8'h18 * io_b_11; // @[ChiselImProc.scala 28:24]
  wire [15:0] _T_35 = _T_32 + _T_33; // @[ChiselImProc.scala 28:13]
  wire [15:0] _T_36 = 8'h24 * io_b_12; // @[ChiselImProc.scala 28:24]
  wire [15:0] _T_38 = _T_35 + _T_36; // @[ChiselImProc.scala 28:13]
  wire [15:0] _T_39 = 8'h18 * io_b_13; // @[ChiselImProc.scala 28:24]
  wire [15:0] _T_41 = _T_38 + _T_39; // @[ChiselImProc.scala 28:13]
  wire [15:0] _T_42 = 8'h6 * io_b_14; // @[ChiselImProc.scala 28:24]
  wire [15:0] _T_44 = _T_41 + _T_42; // @[ChiselImProc.scala 28:13]
  wire [15:0] _T_45 = 8'h4 * io_b_15; // @[ChiselImProc.scala 28:24]
  wire [15:0] _T_47 = _T_44 + _T_45; // @[ChiselImProc.scala 28:13]
  wire [15:0] _T_48 = 8'h10 * io_b_16; // @[ChiselImProc.scala 28:24]
  wire [15:0] _T_50 = _T_47 + _T_48; // @[ChiselImProc.scala 28:13]
  wire [15:0] _T_51 = 8'h18 * io_b_17; // @[ChiselImProc.scala 28:24]
  wire [15:0] _T_53 = _T_50 + _T_51; // @[ChiselImProc.scala 28:13]
  wire [15:0] _T_54 = 8'h10 * io_b_18; // @[ChiselImProc.scala 28:24]
  wire [15:0] _T_56 = _T_53 + _T_54; // @[ChiselImProc.scala 28:13]
  wire [15:0] _T_57 = 8'h4 * io_b_19; // @[ChiselImProc.scala 28:24]
  wire [15:0] _T_59 = _T_56 + _T_57; // @[ChiselImProc.scala 28:13]
  wire [15:0] _T_60 = 8'h1 * io_b_20; // @[ChiselImProc.scala 28:24]
  wire [15:0] _T_62 = _T_59 + _T_60; // @[ChiselImProc.scala 28:13]
  wire [15:0] _T_63 = 8'h4 * io_b_21; // @[ChiselImProc.scala 28:24]
  wire [15:0] _T_65 = _T_62 + _T_63; // @[ChiselImProc.scala 28:13]
  wire [15:0] _T_66 = 8'h6 * io_b_22; // @[ChiselImProc.scala 28:24]
  wire [15:0] _T_68 = _T_65 + _T_66; // @[ChiselImProc.scala 28:13]
  wire [15:0] _T_69 = 8'h4 * io_b_23; // @[ChiselImProc.scala 28:24]
  wire [15:0] _T_71 = _T_68 + _T_69; // @[ChiselImProc.scala 28:13]
  wire [15:0] _T_72 = 8'h1 * io_b_24; // @[ChiselImProc.scala 28:24]
  assign io_output = _T_71 + _T_72; // @[ChiselImProc.scala 31:15]
endmodule
module GaussianBlurFilter(
  input        clock,
  input        reset,
  output       io_enq_ready,
  input        io_enq_valid,
  input  [7:0] io_enq_bits,
  input        io_enq_user,
  input        io_enq_last,
  input        io_deq_ready,
  output       io_deq_valid,
  output [7:0] io_deq_bits,
  output       io_deq_user,
  output       io_deq_last
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
  reg [31:0] _RAND_64;
  reg [31:0] _RAND_65;
  reg [31:0] _RAND_66;
  reg [31:0] _RAND_67;
  reg [31:0] _RAND_68;
  reg [31:0] _RAND_69;
  reg [31:0] _RAND_70;
  reg [31:0] _RAND_71;
  reg [31:0] _RAND_72;
  reg [31:0] _RAND_73;
  reg [31:0] _RAND_74;
  reg [31:0] _RAND_75;
  reg [31:0] _RAND_76;
  reg [31:0] _RAND_77;
  reg [31:0] _RAND_78;
  reg [31:0] _RAND_79;
  reg [31:0] _RAND_80;
  reg [31:0] _RAND_81;
  reg [31:0] _RAND_82;
  reg [31:0] _RAND_83;
  reg [31:0] _RAND_84;
  reg [31:0] _RAND_85;
  reg [31:0] _RAND_86;
  reg [31:0] _RAND_87;
  reg [31:0] _RAND_88;
  reg [31:0] _RAND_89;
  reg [31:0] _RAND_90;
  reg [31:0] _RAND_91;
  reg [31:0] _RAND_92;
  reg [31:0] _RAND_93;
  reg [31:0] _RAND_94;
  reg [31:0] _RAND_95;
  reg [31:0] _RAND_96;
  reg [31:0] _RAND_97;
  reg [31:0] _RAND_98;
  reg [31:0] _RAND_99;
  reg [31:0] _RAND_100;
  reg [31:0] _RAND_101;
  reg [31:0] _RAND_102;
  reg [31:0] _RAND_103;
  reg [31:0] _RAND_104;
  reg [31:0] _RAND_105;
  reg [31:0] _RAND_106;
  reg [31:0] _RAND_107;
  reg [31:0] _RAND_108;
  reg [31:0] _RAND_109;
  reg [31:0] _RAND_110;
  reg [31:0] _RAND_111;
  reg [31:0] _RAND_112;
  reg [31:0] _RAND_113;
  reg [31:0] _RAND_114;
  reg [31:0] _RAND_115;
  reg [31:0] _RAND_116;
  reg [31:0] _RAND_117;
  reg [31:0] _RAND_118;
  reg [31:0] _RAND_119;
  reg [31:0] _RAND_120;
  reg [31:0] _RAND_121;
  reg [31:0] _RAND_122;
  reg [31:0] _RAND_123;
  reg [31:0] _RAND_124;
  reg [31:0] _RAND_125;
  reg [31:0] _RAND_126;
  reg [31:0] _RAND_127;
  reg [31:0] _RAND_128;
  reg [31:0] _RAND_129;
  reg [31:0] _RAND_130;
  reg [31:0] _RAND_131;
  reg [31:0] _RAND_132;
  reg [31:0] _RAND_133;
  reg [31:0] _RAND_134;
  reg [31:0] _RAND_135;
  reg [31:0] _RAND_136;
  reg [31:0] _RAND_137;
  reg [31:0] _RAND_138;
  reg [31:0] _RAND_139;
  reg [31:0] _RAND_140;
  reg [31:0] _RAND_141;
  reg [31:0] _RAND_142;
  reg [31:0] _RAND_143;
  reg [31:0] _RAND_144;
  reg [31:0] _RAND_145;
  reg [31:0] _RAND_146;
  reg [31:0] _RAND_147;
  reg [31:0] _RAND_148;
  reg [31:0] _RAND_149;
  reg [31:0] _RAND_150;
  reg [31:0] _RAND_151;
  reg [31:0] _RAND_152;
  reg [31:0] _RAND_153;
  reg [31:0] _RAND_154;
  reg [31:0] _RAND_155;
  reg [31:0] _RAND_156;
  reg [31:0] _RAND_157;
  reg [31:0] _RAND_158;
  reg [31:0] _RAND_159;
  reg [31:0] _RAND_160;
  reg [31:0] _RAND_161;
  reg [31:0] _RAND_162;
  reg [31:0] _RAND_163;
  reg [31:0] _RAND_164;
  reg [31:0] _RAND_165;
  reg [31:0] _RAND_166;
  reg [31:0] _RAND_167;
  reg [31:0] _RAND_168;
  reg [31:0] _RAND_169;
  reg [31:0] _RAND_170;
  reg [31:0] _RAND_171;
  reg [31:0] _RAND_172;
  reg [31:0] _RAND_173;
  reg [31:0] _RAND_174;
  reg [31:0] _RAND_175;
  reg [31:0] _RAND_176;
  reg [31:0] _RAND_177;
  reg [31:0] _RAND_178;
  reg [31:0] _RAND_179;
  reg [31:0] _RAND_180;
  reg [31:0] _RAND_181;
  reg [31:0] _RAND_182;
  reg [31:0] _RAND_183;
  reg [31:0] _RAND_184;
  reg [31:0] _RAND_185;
  reg [31:0] _RAND_186;
  reg [31:0] _RAND_187;
  reg [31:0] _RAND_188;
  reg [31:0] _RAND_189;
  reg [31:0] _RAND_190;
  reg [31:0] _RAND_191;
  reg [31:0] _RAND_192;
  reg [31:0] _RAND_193;
  reg [31:0] _RAND_194;
  reg [31:0] _RAND_195;
  reg [31:0] _RAND_196;
  reg [31:0] _RAND_197;
  reg [31:0] _RAND_198;
  reg [31:0] _RAND_199;
  reg [31:0] _RAND_200;
  reg [31:0] _RAND_201;
  reg [31:0] _RAND_202;
  reg [31:0] _RAND_203;
  reg [31:0] _RAND_204;
  reg [31:0] _RAND_205;
  reg [31:0] _RAND_206;
  reg [31:0] _RAND_207;
  reg [31:0] _RAND_208;
  reg [31:0] _RAND_209;
  reg [31:0] _RAND_210;
  reg [31:0] _RAND_211;
  reg [31:0] _RAND_212;
  reg [31:0] _RAND_213;
  reg [31:0] _RAND_214;
  reg [31:0] _RAND_215;
  reg [31:0] _RAND_216;
  reg [31:0] _RAND_217;
  reg [31:0] _RAND_218;
  reg [31:0] _RAND_219;
  reg [31:0] _RAND_220;
  reg [31:0] _RAND_221;
  reg [31:0] _RAND_222;
  reg [31:0] _RAND_223;
  reg [31:0] _RAND_224;
  reg [31:0] _RAND_225;
  reg [31:0] _RAND_226;
  reg [31:0] _RAND_227;
  reg [31:0] _RAND_228;
  reg [31:0] _RAND_229;
  reg [31:0] _RAND_230;
  reg [31:0] _RAND_231;
  reg [31:0] _RAND_232;
  reg [31:0] _RAND_233;
  reg [31:0] _RAND_234;
  reg [31:0] _RAND_235;
  reg [31:0] _RAND_236;
  reg [31:0] _RAND_237;
  reg [31:0] _RAND_238;
  reg [31:0] _RAND_239;
  reg [31:0] _RAND_240;
  reg [31:0] _RAND_241;
  reg [31:0] _RAND_242;
  reg [31:0] _RAND_243;
  reg [31:0] _RAND_244;
  reg [31:0] _RAND_245;
  reg [31:0] _RAND_246;
  reg [31:0] _RAND_247;
  reg [31:0] _RAND_248;
  reg [31:0] _RAND_249;
  reg [31:0] _RAND_250;
  reg [31:0] _RAND_251;
  reg [31:0] _RAND_252;
  reg [31:0] _RAND_253;
  reg [31:0] _RAND_254;
  reg [31:0] _RAND_255;
  reg [31:0] _RAND_256;
  reg [31:0] _RAND_257;
  reg [31:0] _RAND_258;
  reg [31:0] _RAND_259;
  reg [31:0] _RAND_260;
  reg [31:0] _RAND_261;
  reg [31:0] _RAND_262;
  reg [31:0] _RAND_263;
  reg [31:0] _RAND_264;
  reg [31:0] _RAND_265;
  reg [31:0] _RAND_266;
  reg [31:0] _RAND_267;
  reg [31:0] _RAND_268;
  reg [31:0] _RAND_269;
  reg [31:0] _RAND_270;
  reg [31:0] _RAND_271;
  reg [31:0] _RAND_272;
  reg [31:0] _RAND_273;
  reg [31:0] _RAND_274;
  reg [31:0] _RAND_275;
  reg [31:0] _RAND_276;
  reg [31:0] _RAND_277;
  reg [31:0] _RAND_278;
  reg [31:0] _RAND_279;
  reg [31:0] _RAND_280;
  reg [31:0] _RAND_281;
  reg [31:0] _RAND_282;
  reg [31:0] _RAND_283;
  reg [31:0] _RAND_284;
  reg [31:0] _RAND_285;
  reg [31:0] _RAND_286;
  reg [31:0] _RAND_287;
  reg [31:0] _RAND_288;
  reg [31:0] _RAND_289;
  reg [31:0] _RAND_290;
  reg [31:0] _RAND_291;
  reg [31:0] _RAND_292;
  reg [31:0] _RAND_293;
  reg [31:0] _RAND_294;
  reg [31:0] _RAND_295;
  reg [31:0] _RAND_296;
  reg [31:0] _RAND_297;
  reg [31:0] _RAND_298;
  reg [31:0] _RAND_299;
  reg [31:0] _RAND_300;
  reg [31:0] _RAND_301;
  reg [31:0] _RAND_302;
  reg [31:0] _RAND_303;
  reg [31:0] _RAND_304;
  reg [31:0] _RAND_305;
  reg [31:0] _RAND_306;
  reg [31:0] _RAND_307;
  reg [31:0] _RAND_308;
  reg [31:0] _RAND_309;
  reg [31:0] _RAND_310;
  reg [31:0] _RAND_311;
  reg [31:0] _RAND_312;
  reg [31:0] _RAND_313;
  reg [31:0] _RAND_314;
  reg [31:0] _RAND_315;
  reg [31:0] _RAND_316;
  reg [31:0] _RAND_317;
  reg [31:0] _RAND_318;
  reg [31:0] _RAND_319;
  reg [31:0] _RAND_320;
  reg [31:0] _RAND_321;
  reg [31:0] _RAND_322;
  reg [31:0] _RAND_323;
  reg [31:0] _RAND_324;
  reg [31:0] _RAND_325;
  reg [31:0] _RAND_326;
  reg [31:0] _RAND_327;
  reg [31:0] _RAND_328;
  reg [31:0] _RAND_329;
  reg [31:0] _RAND_330;
  reg [31:0] _RAND_331;
  reg [31:0] _RAND_332;
  reg [31:0] _RAND_333;
  reg [31:0] _RAND_334;
  reg [31:0] _RAND_335;
  reg [31:0] _RAND_336;
  reg [31:0] _RAND_337;
  reg [31:0] _RAND_338;
  reg [31:0] _RAND_339;
  reg [31:0] _RAND_340;
  reg [31:0] _RAND_341;
  reg [31:0] _RAND_342;
  reg [31:0] _RAND_343;
  reg [31:0] _RAND_344;
  reg [31:0] _RAND_345;
  reg [31:0] _RAND_346;
  reg [31:0] _RAND_347;
  reg [31:0] _RAND_348;
  reg [31:0] _RAND_349;
  reg [31:0] _RAND_350;
  reg [31:0] _RAND_351;
  reg [31:0] _RAND_352;
  reg [31:0] _RAND_353;
  reg [31:0] _RAND_354;
  reg [31:0] _RAND_355;
  reg [31:0] _RAND_356;
  reg [31:0] _RAND_357;
  reg [31:0] _RAND_358;
  reg [31:0] _RAND_359;
  reg [31:0] _RAND_360;
  reg [31:0] _RAND_361;
  reg [31:0] _RAND_362;
  reg [31:0] _RAND_363;
  reg [31:0] _RAND_364;
  reg [31:0] _RAND_365;
  reg [31:0] _RAND_366;
  reg [31:0] _RAND_367;
  reg [31:0] _RAND_368;
  reg [31:0] _RAND_369;
  reg [31:0] _RAND_370;
  reg [31:0] _RAND_371;
  reg [31:0] _RAND_372;
  reg [31:0] _RAND_373;
  reg [31:0] _RAND_374;
  reg [31:0] _RAND_375;
  reg [31:0] _RAND_376;
  reg [31:0] _RAND_377;
  reg [31:0] _RAND_378;
  reg [31:0] _RAND_379;
  reg [31:0] _RAND_380;
  reg [31:0] _RAND_381;
  reg [31:0] _RAND_382;
  reg [31:0] _RAND_383;
  reg [31:0] _RAND_384;
  reg [31:0] _RAND_385;
  reg [31:0] _RAND_386;
  reg [31:0] _RAND_387;
  reg [31:0] _RAND_388;
  reg [31:0] _RAND_389;
  reg [31:0] _RAND_390;
  reg [31:0] _RAND_391;
  reg [31:0] _RAND_392;
  reg [31:0] _RAND_393;
  reg [31:0] _RAND_394;
  reg [31:0] _RAND_395;
  reg [31:0] _RAND_396;
  reg [31:0] _RAND_397;
  reg [31:0] _RAND_398;
  reg [31:0] _RAND_399;
  reg [31:0] _RAND_400;
  reg [31:0] _RAND_401;
  reg [31:0] _RAND_402;
  reg [31:0] _RAND_403;
  reg [31:0] _RAND_404;
  reg [31:0] _RAND_405;
  reg [31:0] _RAND_406;
  reg [31:0] _RAND_407;
  reg [31:0] _RAND_408;
  reg [31:0] _RAND_409;
  reg [31:0] _RAND_410;
  reg [31:0] _RAND_411;
  reg [31:0] _RAND_412;
  reg [31:0] _RAND_413;
  reg [31:0] _RAND_414;
  reg [31:0] _RAND_415;
  reg [31:0] _RAND_416;
  reg [31:0] _RAND_417;
  reg [31:0] _RAND_418;
  reg [31:0] _RAND_419;
  reg [31:0] _RAND_420;
  reg [31:0] _RAND_421;
  reg [31:0] _RAND_422;
  reg [31:0] _RAND_423;
  reg [31:0] _RAND_424;
  reg [31:0] _RAND_425;
  reg [31:0] _RAND_426;
  reg [31:0] _RAND_427;
  reg [31:0] _RAND_428;
  reg [31:0] _RAND_429;
  reg [31:0] _RAND_430;
  reg [31:0] _RAND_431;
  reg [31:0] _RAND_432;
  reg [31:0] _RAND_433;
  reg [31:0] _RAND_434;
  reg [31:0] _RAND_435;
  reg [31:0] _RAND_436;
  reg [31:0] _RAND_437;
  reg [31:0] _RAND_438;
  reg [31:0] _RAND_439;
  reg [31:0] _RAND_440;
  reg [31:0] _RAND_441;
  reg [31:0] _RAND_442;
  reg [31:0] _RAND_443;
  reg [31:0] _RAND_444;
  reg [31:0] _RAND_445;
  reg [31:0] _RAND_446;
  reg [31:0] _RAND_447;
  reg [31:0] _RAND_448;
  reg [31:0] _RAND_449;
  reg [31:0] _RAND_450;
  reg [31:0] _RAND_451;
  reg [31:0] _RAND_452;
  reg [31:0] _RAND_453;
  reg [31:0] _RAND_454;
  reg [31:0] _RAND_455;
  reg [31:0] _RAND_456;
  reg [31:0] _RAND_457;
  reg [31:0] _RAND_458;
  reg [31:0] _RAND_459;
  reg [31:0] _RAND_460;
  reg [31:0] _RAND_461;
  reg [31:0] _RAND_462;
  reg [31:0] _RAND_463;
  reg [31:0] _RAND_464;
  reg [31:0] _RAND_465;
  reg [31:0] _RAND_466;
  reg [31:0] _RAND_467;
  reg [31:0] _RAND_468;
  reg [31:0] _RAND_469;
  reg [31:0] _RAND_470;
  reg [31:0] _RAND_471;
  reg [31:0] _RAND_472;
  reg [31:0] _RAND_473;
  reg [31:0] _RAND_474;
  reg [31:0] _RAND_475;
  reg [31:0] _RAND_476;
  reg [31:0] _RAND_477;
  reg [31:0] _RAND_478;
  reg [31:0] _RAND_479;
  reg [31:0] _RAND_480;
  reg [31:0] _RAND_481;
  reg [31:0] _RAND_482;
  reg [31:0] _RAND_483;
  reg [31:0] _RAND_484;
  reg [31:0] _RAND_485;
  reg [31:0] _RAND_486;
  reg [31:0] _RAND_487;
  reg [31:0] _RAND_488;
  reg [31:0] _RAND_489;
  reg [31:0] _RAND_490;
  reg [31:0] _RAND_491;
  reg [31:0] _RAND_492;
  reg [31:0] _RAND_493;
  reg [31:0] _RAND_494;
  reg [31:0] _RAND_495;
  reg [31:0] _RAND_496;
  reg [31:0] _RAND_497;
  reg [31:0] _RAND_498;
  reg [31:0] _RAND_499;
  reg [31:0] _RAND_500;
  reg [31:0] _RAND_501;
  reg [31:0] _RAND_502;
  reg [31:0] _RAND_503;
  reg [31:0] _RAND_504;
  reg [31:0] _RAND_505;
  reg [31:0] _RAND_506;
  reg [31:0] _RAND_507;
  reg [31:0] _RAND_508;
  reg [31:0] _RAND_509;
  reg [31:0] _RAND_510;
  reg [31:0] _RAND_511;
  reg [31:0] _RAND_512;
  reg [31:0] _RAND_513;
  reg [31:0] _RAND_514;
  reg [31:0] _RAND_515;
  reg [31:0] _RAND_516;
  reg [31:0] _RAND_517;
  reg [31:0] _RAND_518;
  reg [31:0] _RAND_519;
  reg [31:0] _RAND_520;
  reg [31:0] _RAND_521;
  reg [31:0] _RAND_522;
  reg [31:0] _RAND_523;
  reg [31:0] _RAND_524;
  reg [31:0] _RAND_525;
  reg [31:0] _RAND_526;
  reg [31:0] _RAND_527;
  reg [31:0] _RAND_528;
  reg [31:0] _RAND_529;
  reg [31:0] _RAND_530;
  reg [31:0] _RAND_531;
  reg [31:0] _RAND_532;
  reg [31:0] _RAND_533;
  reg [31:0] _RAND_534;
  reg [31:0] _RAND_535;
  reg [31:0] _RAND_536;
  reg [31:0] _RAND_537;
  reg [31:0] _RAND_538;
  reg [31:0] _RAND_539;
  reg [31:0] _RAND_540;
  reg [31:0] _RAND_541;
  reg [31:0] _RAND_542;
  reg [31:0] _RAND_543;
  reg [31:0] _RAND_544;
  reg [31:0] _RAND_545;
  reg [31:0] _RAND_546;
  reg [31:0] _RAND_547;
  reg [31:0] _RAND_548;
  reg [31:0] _RAND_549;
  reg [31:0] _RAND_550;
  reg [31:0] _RAND_551;
  reg [31:0] _RAND_552;
  reg [31:0] _RAND_553;
  reg [31:0] _RAND_554;
  reg [31:0] _RAND_555;
  reg [31:0] _RAND_556;
  reg [31:0] _RAND_557;
  reg [31:0] _RAND_558;
  reg [31:0] _RAND_559;
  reg [31:0] _RAND_560;
  reg [31:0] _RAND_561;
  reg [31:0] _RAND_562;
  reg [31:0] _RAND_563;
  reg [31:0] _RAND_564;
  reg [31:0] _RAND_565;
  reg [31:0] _RAND_566;
  reg [31:0] _RAND_567;
  reg [31:0] _RAND_568;
  reg [31:0] _RAND_569;
  reg [31:0] _RAND_570;
  reg [31:0] _RAND_571;
  reg [31:0] _RAND_572;
  reg [31:0] _RAND_573;
  reg [31:0] _RAND_574;
  reg [31:0] _RAND_575;
  reg [31:0] _RAND_576;
  reg [31:0] _RAND_577;
  reg [31:0] _RAND_578;
  reg [31:0] _RAND_579;
  reg [31:0] _RAND_580;
  reg [31:0] _RAND_581;
  reg [31:0] _RAND_582;
  reg [31:0] _RAND_583;
  reg [31:0] _RAND_584;
  reg [31:0] _RAND_585;
  reg [31:0] _RAND_586;
  reg [31:0] _RAND_587;
  reg [31:0] _RAND_588;
  reg [31:0] _RAND_589;
  reg [31:0] _RAND_590;
  reg [31:0] _RAND_591;
  reg [31:0] _RAND_592;
  reg [31:0] _RAND_593;
  reg [31:0] _RAND_594;
  reg [31:0] _RAND_595;
  reg [31:0] _RAND_596;
  reg [31:0] _RAND_597;
  reg [31:0] _RAND_598;
  reg [31:0] _RAND_599;
  reg [31:0] _RAND_600;
  reg [31:0] _RAND_601;
  reg [31:0] _RAND_602;
  reg [31:0] _RAND_603;
  reg [31:0] _RAND_604;
  reg [31:0] _RAND_605;
  reg [31:0] _RAND_606;
  reg [31:0] _RAND_607;
  reg [31:0] _RAND_608;
  reg [31:0] _RAND_609;
  reg [31:0] _RAND_610;
  reg [31:0] _RAND_611;
  reg [31:0] _RAND_612;
  reg [31:0] _RAND_613;
  reg [31:0] _RAND_614;
  reg [31:0] _RAND_615;
  reg [31:0] _RAND_616;
  reg [31:0] _RAND_617;
  reg [31:0] _RAND_618;
  reg [31:0] _RAND_619;
  reg [31:0] _RAND_620;
  reg [31:0] _RAND_621;
  reg [31:0] _RAND_622;
  reg [31:0] _RAND_623;
  reg [31:0] _RAND_624;
  reg [31:0] _RAND_625;
  reg [31:0] _RAND_626;
  reg [31:0] _RAND_627;
  reg [31:0] _RAND_628;
  reg [31:0] _RAND_629;
  reg [31:0] _RAND_630;
  reg [31:0] _RAND_631;
  reg [31:0] _RAND_632;
  reg [31:0] _RAND_633;
  reg [31:0] _RAND_634;
  reg [31:0] _RAND_635;
  reg [31:0] _RAND_636;
  reg [31:0] _RAND_637;
  reg [31:0] _RAND_638;
  reg [31:0] _RAND_639;
  reg [31:0] _RAND_640;
  reg [31:0] _RAND_641;
  reg [31:0] _RAND_642;
  reg [31:0] _RAND_643;
  reg [31:0] _RAND_644;
  reg [31:0] _RAND_645;
  reg [31:0] _RAND_646;
  reg [31:0] _RAND_647;
  reg [31:0] _RAND_648;
  reg [31:0] _RAND_649;
  reg [31:0] _RAND_650;
  reg [31:0] _RAND_651;
  reg [31:0] _RAND_652;
  reg [31:0] _RAND_653;
  reg [31:0] _RAND_654;
  reg [31:0] _RAND_655;
  reg [31:0] _RAND_656;
  reg [31:0] _RAND_657;
  reg [31:0] _RAND_658;
  reg [31:0] _RAND_659;
  reg [31:0] _RAND_660;
  reg [31:0] _RAND_661;
  reg [31:0] _RAND_662;
  reg [31:0] _RAND_663;
  reg [31:0] _RAND_664;
  reg [31:0] _RAND_665;
  reg [31:0] _RAND_666;
  reg [31:0] _RAND_667;
  reg [31:0] _RAND_668;
  reg [31:0] _RAND_669;
  reg [31:0] _RAND_670;
  reg [31:0] _RAND_671;
  reg [31:0] _RAND_672;
  reg [31:0] _RAND_673;
  reg [31:0] _RAND_674;
  reg [31:0] _RAND_675;
  reg [31:0] _RAND_676;
  reg [31:0] _RAND_677;
  reg [31:0] _RAND_678;
  reg [31:0] _RAND_679;
  reg [31:0] _RAND_680;
  reg [31:0] _RAND_681;
  reg [31:0] _RAND_682;
  reg [31:0] _RAND_683;
  reg [31:0] _RAND_684;
  reg [31:0] _RAND_685;
  reg [31:0] _RAND_686;
  reg [31:0] _RAND_687;
  reg [31:0] _RAND_688;
  reg [31:0] _RAND_689;
  reg [31:0] _RAND_690;
  reg [31:0] _RAND_691;
  reg [31:0] _RAND_692;
  reg [31:0] _RAND_693;
  reg [31:0] _RAND_694;
  reg [31:0] _RAND_695;
  reg [31:0] _RAND_696;
  reg [31:0] _RAND_697;
  reg [31:0] _RAND_698;
  reg [31:0] _RAND_699;
  reg [31:0] _RAND_700;
  reg [31:0] _RAND_701;
  reg [31:0] _RAND_702;
  reg [31:0] _RAND_703;
  reg [31:0] _RAND_704;
  reg [31:0] _RAND_705;
  reg [31:0] _RAND_706;
  reg [31:0] _RAND_707;
  reg [31:0] _RAND_708;
  reg [31:0] _RAND_709;
  reg [31:0] _RAND_710;
  reg [31:0] _RAND_711;
  reg [31:0] _RAND_712;
  reg [31:0] _RAND_713;
  reg [31:0] _RAND_714;
  reg [31:0] _RAND_715;
  reg [31:0] _RAND_716;
  reg [31:0] _RAND_717;
  reg [31:0] _RAND_718;
  reg [31:0] _RAND_719;
  reg [31:0] _RAND_720;
  reg [31:0] _RAND_721;
  reg [31:0] _RAND_722;
  reg [31:0] _RAND_723;
  reg [31:0] _RAND_724;
  reg [31:0] _RAND_725;
  reg [31:0] _RAND_726;
  reg [31:0] _RAND_727;
  reg [31:0] _RAND_728;
  reg [31:0] _RAND_729;
  reg [31:0] _RAND_730;
  reg [31:0] _RAND_731;
  reg [31:0] _RAND_732;
  reg [31:0] _RAND_733;
  reg [31:0] _RAND_734;
  reg [31:0] _RAND_735;
  reg [31:0] _RAND_736;
  reg [31:0] _RAND_737;
  reg [31:0] _RAND_738;
  reg [31:0] _RAND_739;
  reg [31:0] _RAND_740;
  reg [31:0] _RAND_741;
  reg [31:0] _RAND_742;
  reg [31:0] _RAND_743;
  reg [31:0] _RAND_744;
  reg [31:0] _RAND_745;
  reg [31:0] _RAND_746;
  reg [31:0] _RAND_747;
  reg [31:0] _RAND_748;
  reg [31:0] _RAND_749;
  reg [31:0] _RAND_750;
  reg [31:0] _RAND_751;
  reg [31:0] _RAND_752;
  reg [31:0] _RAND_753;
  reg [31:0] _RAND_754;
  reg [31:0] _RAND_755;
  reg [31:0] _RAND_756;
  reg [31:0] _RAND_757;
  reg [31:0] _RAND_758;
  reg [31:0] _RAND_759;
  reg [31:0] _RAND_760;
  reg [31:0] _RAND_761;
  reg [31:0] _RAND_762;
  reg [31:0] _RAND_763;
  reg [31:0] _RAND_764;
  reg [31:0] _RAND_765;
  reg [31:0] _RAND_766;
  reg [31:0] _RAND_767;
  reg [31:0] _RAND_768;
  reg [31:0] _RAND_769;
  reg [31:0] _RAND_770;
  reg [31:0] _RAND_771;
  reg [31:0] _RAND_772;
  reg [31:0] _RAND_773;
  reg [31:0] _RAND_774;
  reg [31:0] _RAND_775;
  reg [31:0] _RAND_776;
  reg [31:0] _RAND_777;
  reg [31:0] _RAND_778;
  reg [31:0] _RAND_779;
  reg [31:0] _RAND_780;
  reg [31:0] _RAND_781;
  reg [31:0] _RAND_782;
  reg [31:0] _RAND_783;
  reg [31:0] _RAND_784;
  reg [31:0] _RAND_785;
  reg [31:0] _RAND_786;
  reg [31:0] _RAND_787;
  reg [31:0] _RAND_788;
  reg [31:0] _RAND_789;
  reg [31:0] _RAND_790;
  reg [31:0] _RAND_791;
  reg [31:0] _RAND_792;
  reg [31:0] _RAND_793;
  reg [31:0] _RAND_794;
  reg [31:0] _RAND_795;
  reg [31:0] _RAND_796;
  reg [31:0] _RAND_797;
  reg [31:0] _RAND_798;
  reg [31:0] _RAND_799;
  reg [31:0] _RAND_800;
  reg [31:0] _RAND_801;
  reg [31:0] _RAND_802;
  reg [31:0] _RAND_803;
  reg [31:0] _RAND_804;
  reg [31:0] _RAND_805;
  reg [31:0] _RAND_806;
  reg [31:0] _RAND_807;
  reg [31:0] _RAND_808;
  reg [31:0] _RAND_809;
  reg [31:0] _RAND_810;
  reg [31:0] _RAND_811;
  reg [31:0] _RAND_812;
  reg [31:0] _RAND_813;
  reg [31:0] _RAND_814;
  reg [31:0] _RAND_815;
  reg [31:0] _RAND_816;
  reg [31:0] _RAND_817;
  reg [31:0] _RAND_818;
  reg [31:0] _RAND_819;
  reg [31:0] _RAND_820;
  reg [31:0] _RAND_821;
  reg [31:0] _RAND_822;
  reg [31:0] _RAND_823;
  reg [31:0] _RAND_824;
  reg [31:0] _RAND_825;
  reg [31:0] _RAND_826;
  reg [31:0] _RAND_827;
  reg [31:0] _RAND_828;
  reg [31:0] _RAND_829;
  reg [31:0] _RAND_830;
  reg [31:0] _RAND_831;
  reg [31:0] _RAND_832;
  reg [31:0] _RAND_833;
  reg [31:0] _RAND_834;
  reg [31:0] _RAND_835;
  reg [31:0] _RAND_836;
  reg [31:0] _RAND_837;
  reg [31:0] _RAND_838;
  reg [31:0] _RAND_839;
  reg [31:0] _RAND_840;
  reg [31:0] _RAND_841;
  reg [31:0] _RAND_842;
  reg [31:0] _RAND_843;
  reg [31:0] _RAND_844;
  reg [31:0] _RAND_845;
  reg [31:0] _RAND_846;
  reg [31:0] _RAND_847;
  reg [31:0] _RAND_848;
  reg [31:0] _RAND_849;
  reg [31:0] _RAND_850;
  reg [31:0] _RAND_851;
  reg [31:0] _RAND_852;
  reg [31:0] _RAND_853;
  reg [31:0] _RAND_854;
  reg [31:0] _RAND_855;
  reg [31:0] _RAND_856;
  reg [31:0] _RAND_857;
  reg [31:0] _RAND_858;
  reg [31:0] _RAND_859;
  reg [31:0] _RAND_860;
  reg [31:0] _RAND_861;
  reg [31:0] _RAND_862;
  reg [31:0] _RAND_863;
  reg [31:0] _RAND_864;
  reg [31:0] _RAND_865;
  reg [31:0] _RAND_866;
  reg [31:0] _RAND_867;
  reg [31:0] _RAND_868;
  reg [31:0] _RAND_869;
  reg [31:0] _RAND_870;
  reg [31:0] _RAND_871;
  reg [31:0] _RAND_872;
  reg [31:0] _RAND_873;
  reg [31:0] _RAND_874;
  reg [31:0] _RAND_875;
  reg [31:0] _RAND_876;
  reg [31:0] _RAND_877;
  reg [31:0] _RAND_878;
  reg [31:0] _RAND_879;
  reg [31:0] _RAND_880;
  reg [31:0] _RAND_881;
  reg [31:0] _RAND_882;
  reg [31:0] _RAND_883;
  reg [31:0] _RAND_884;
  reg [31:0] _RAND_885;
  reg [31:0] _RAND_886;
  reg [31:0] _RAND_887;
  reg [31:0] _RAND_888;
  reg [31:0] _RAND_889;
  reg [31:0] _RAND_890;
  reg [31:0] _RAND_891;
  reg [31:0] _RAND_892;
  reg [31:0] _RAND_893;
  reg [31:0] _RAND_894;
  reg [31:0] _RAND_895;
  reg [31:0] _RAND_896;
  reg [31:0] _RAND_897;
  reg [31:0] _RAND_898;
  reg [31:0] _RAND_899;
  reg [31:0] _RAND_900;
  reg [31:0] _RAND_901;
  reg [31:0] _RAND_902;
  reg [31:0] _RAND_903;
  reg [31:0] _RAND_904;
  reg [31:0] _RAND_905;
  reg [31:0] _RAND_906;
  reg [31:0] _RAND_907;
  reg [31:0] _RAND_908;
  reg [31:0] _RAND_909;
  reg [31:0] _RAND_910;
  reg [31:0] _RAND_911;
  reg [31:0] _RAND_912;
  reg [31:0] _RAND_913;
  reg [31:0] _RAND_914;
  reg [31:0] _RAND_915;
  reg [31:0] _RAND_916;
  reg [31:0] _RAND_917;
  reg [31:0] _RAND_918;
  reg [31:0] _RAND_919;
  reg [31:0] _RAND_920;
  reg [31:0] _RAND_921;
  reg [31:0] _RAND_922;
  reg [31:0] _RAND_923;
  reg [31:0] _RAND_924;
  reg [31:0] _RAND_925;
  reg [31:0] _RAND_926;
  reg [31:0] _RAND_927;
  reg [31:0] _RAND_928;
  reg [31:0] _RAND_929;
  reg [31:0] _RAND_930;
  reg [31:0] _RAND_931;
  reg [31:0] _RAND_932;
  reg [31:0] _RAND_933;
  reg [31:0] _RAND_934;
  reg [31:0] _RAND_935;
  reg [31:0] _RAND_936;
  reg [31:0] _RAND_937;
  reg [31:0] _RAND_938;
  reg [31:0] _RAND_939;
  reg [31:0] _RAND_940;
  reg [31:0] _RAND_941;
  reg [31:0] _RAND_942;
  reg [31:0] _RAND_943;
  reg [31:0] _RAND_944;
  reg [31:0] _RAND_945;
  reg [31:0] _RAND_946;
  reg [31:0] _RAND_947;
  reg [31:0] _RAND_948;
  reg [31:0] _RAND_949;
  reg [31:0] _RAND_950;
  reg [31:0] _RAND_951;
  reg [31:0] _RAND_952;
  reg [31:0] _RAND_953;
  reg [31:0] _RAND_954;
  reg [31:0] _RAND_955;
  reg [31:0] _RAND_956;
  reg [31:0] _RAND_957;
  reg [31:0] _RAND_958;
  reg [31:0] _RAND_959;
  reg [31:0] _RAND_960;
  reg [31:0] _RAND_961;
  reg [31:0] _RAND_962;
  reg [31:0] _RAND_963;
  reg [31:0] _RAND_964;
  reg [31:0] _RAND_965;
  reg [31:0] _RAND_966;
  reg [31:0] _RAND_967;
  reg [31:0] _RAND_968;
  reg [31:0] _RAND_969;
  reg [31:0] _RAND_970;
  reg [31:0] _RAND_971;
  reg [31:0] _RAND_972;
  reg [31:0] _RAND_973;
  reg [31:0] _RAND_974;
  reg [31:0] _RAND_975;
  reg [31:0] _RAND_976;
  reg [31:0] _RAND_977;
  reg [31:0] _RAND_978;
  reg [31:0] _RAND_979;
  reg [31:0] _RAND_980;
  reg [31:0] _RAND_981;
  reg [31:0] _RAND_982;
  reg [31:0] _RAND_983;
  reg [31:0] _RAND_984;
  reg [31:0] _RAND_985;
  reg [31:0] _RAND_986;
  reg [31:0] _RAND_987;
  reg [31:0] _RAND_988;
  reg [31:0] _RAND_989;
  reg [31:0] _RAND_990;
  reg [31:0] _RAND_991;
  reg [31:0] _RAND_992;
  reg [31:0] _RAND_993;
  reg [31:0] _RAND_994;
  reg [31:0] _RAND_995;
  reg [31:0] _RAND_996;
  reg [31:0] _RAND_997;
  reg [31:0] _RAND_998;
  reg [31:0] _RAND_999;
  reg [31:0] _RAND_1000;
  reg [31:0] _RAND_1001;
  reg [31:0] _RAND_1002;
  reg [31:0] _RAND_1003;
  reg [31:0] _RAND_1004;
  reg [31:0] _RAND_1005;
  reg [31:0] _RAND_1006;
  reg [31:0] _RAND_1007;
  reg [31:0] _RAND_1008;
  reg [31:0] _RAND_1009;
  reg [31:0] _RAND_1010;
  reg [31:0] _RAND_1011;
  reg [31:0] _RAND_1012;
  reg [31:0] _RAND_1013;
  reg [31:0] _RAND_1014;
  reg [31:0] _RAND_1015;
  reg [31:0] _RAND_1016;
  reg [31:0] _RAND_1017;
  reg [31:0] _RAND_1018;
  reg [31:0] _RAND_1019;
  reg [31:0] _RAND_1020;
  reg [31:0] _RAND_1021;
  reg [31:0] _RAND_1022;
  reg [31:0] _RAND_1023;
  reg [31:0] _RAND_1024;
  reg [31:0] _RAND_1025;
  reg [31:0] _RAND_1026;
  reg [31:0] _RAND_1027;
  reg [31:0] _RAND_1028;
  reg [31:0] _RAND_1029;
  reg [31:0] _RAND_1030;
  reg [31:0] _RAND_1031;
  reg [31:0] _RAND_1032;
  reg [31:0] _RAND_1033;
  reg [31:0] _RAND_1034;
  reg [31:0] _RAND_1035;
  reg [31:0] _RAND_1036;
  reg [31:0] _RAND_1037;
  reg [31:0] _RAND_1038;
  reg [31:0] _RAND_1039;
  reg [31:0] _RAND_1040;
  reg [31:0] _RAND_1041;
  reg [31:0] _RAND_1042;
  reg [31:0] _RAND_1043;
  reg [31:0] _RAND_1044;
  reg [31:0] _RAND_1045;
  reg [31:0] _RAND_1046;
  reg [31:0] _RAND_1047;
  reg [31:0] _RAND_1048;
  reg [31:0] _RAND_1049;
  reg [31:0] _RAND_1050;
  reg [31:0] _RAND_1051;
  reg [31:0] _RAND_1052;
  reg [31:0] _RAND_1053;
  reg [31:0] _RAND_1054;
  reg [31:0] _RAND_1055;
  reg [31:0] _RAND_1056;
  reg [31:0] _RAND_1057;
  reg [31:0] _RAND_1058;
  reg [31:0] _RAND_1059;
  reg [31:0] _RAND_1060;
  reg [31:0] _RAND_1061;
  reg [31:0] _RAND_1062;
  reg [31:0] _RAND_1063;
  reg [31:0] _RAND_1064;
  reg [31:0] _RAND_1065;
  reg [31:0] _RAND_1066;
  reg [31:0] _RAND_1067;
  reg [31:0] _RAND_1068;
  reg [31:0] _RAND_1069;
  reg [31:0] _RAND_1070;
  reg [31:0] _RAND_1071;
  reg [31:0] _RAND_1072;
  reg [31:0] _RAND_1073;
  reg [31:0] _RAND_1074;
  reg [31:0] _RAND_1075;
  reg [31:0] _RAND_1076;
  reg [31:0] _RAND_1077;
  reg [31:0] _RAND_1078;
  reg [31:0] _RAND_1079;
  reg [31:0] _RAND_1080;
  reg [31:0] _RAND_1081;
  reg [31:0] _RAND_1082;
  reg [31:0] _RAND_1083;
  reg [31:0] _RAND_1084;
  reg [31:0] _RAND_1085;
  reg [31:0] _RAND_1086;
  reg [31:0] _RAND_1087;
  reg [31:0] _RAND_1088;
  reg [31:0] _RAND_1089;
  reg [31:0] _RAND_1090;
  reg [31:0] _RAND_1091;
  reg [31:0] _RAND_1092;
  reg [31:0] _RAND_1093;
  reg [31:0] _RAND_1094;
  reg [31:0] _RAND_1095;
  reg [31:0] _RAND_1096;
  reg [31:0] _RAND_1097;
  reg [31:0] _RAND_1098;
  reg [31:0] _RAND_1099;
  reg [31:0] _RAND_1100;
  reg [31:0] _RAND_1101;
  reg [31:0] _RAND_1102;
  reg [31:0] _RAND_1103;
  reg [31:0] _RAND_1104;
  reg [31:0] _RAND_1105;
  reg [31:0] _RAND_1106;
  reg [31:0] _RAND_1107;
  reg [31:0] _RAND_1108;
  reg [31:0] _RAND_1109;
  reg [31:0] _RAND_1110;
  reg [31:0] _RAND_1111;
  reg [31:0] _RAND_1112;
  reg [31:0] _RAND_1113;
  reg [31:0] _RAND_1114;
  reg [31:0] _RAND_1115;
  reg [31:0] _RAND_1116;
  reg [31:0] _RAND_1117;
  reg [31:0] _RAND_1118;
  reg [31:0] _RAND_1119;
  reg [31:0] _RAND_1120;
  reg [31:0] _RAND_1121;
  reg [31:0] _RAND_1122;
  reg [31:0] _RAND_1123;
  reg [31:0] _RAND_1124;
  reg [31:0] _RAND_1125;
  reg [31:0] _RAND_1126;
  reg [31:0] _RAND_1127;
  reg [31:0] _RAND_1128;
  reg [31:0] _RAND_1129;
  reg [31:0] _RAND_1130;
  reg [31:0] _RAND_1131;
  reg [31:0] _RAND_1132;
  reg [31:0] _RAND_1133;
  reg [31:0] _RAND_1134;
  reg [31:0] _RAND_1135;
  reg [31:0] _RAND_1136;
  reg [31:0] _RAND_1137;
  reg [31:0] _RAND_1138;
  reg [31:0] _RAND_1139;
  reg [31:0] _RAND_1140;
  reg [31:0] _RAND_1141;
  reg [31:0] _RAND_1142;
  reg [31:0] _RAND_1143;
  reg [31:0] _RAND_1144;
  reg [31:0] _RAND_1145;
  reg [31:0] _RAND_1146;
  reg [31:0] _RAND_1147;
  reg [31:0] _RAND_1148;
  reg [31:0] _RAND_1149;
  reg [31:0] _RAND_1150;
  reg [31:0] _RAND_1151;
  reg [31:0] _RAND_1152;
  reg [31:0] _RAND_1153;
  reg [31:0] _RAND_1154;
  reg [31:0] _RAND_1155;
  reg [31:0] _RAND_1156;
  reg [31:0] _RAND_1157;
  reg [31:0] _RAND_1158;
  reg [31:0] _RAND_1159;
  reg [31:0] _RAND_1160;
  reg [31:0] _RAND_1161;
  reg [31:0] _RAND_1162;
  reg [31:0] _RAND_1163;
  reg [31:0] _RAND_1164;
  reg [31:0] _RAND_1165;
  reg [31:0] _RAND_1166;
  reg [31:0] _RAND_1167;
  reg [31:0] _RAND_1168;
  reg [31:0] _RAND_1169;
  reg [31:0] _RAND_1170;
  reg [31:0] _RAND_1171;
  reg [31:0] _RAND_1172;
  reg [31:0] _RAND_1173;
  reg [31:0] _RAND_1174;
  reg [31:0] _RAND_1175;
  reg [31:0] _RAND_1176;
  reg [31:0] _RAND_1177;
  reg [31:0] _RAND_1178;
  reg [31:0] _RAND_1179;
  reg [31:0] _RAND_1180;
  reg [31:0] _RAND_1181;
  reg [31:0] _RAND_1182;
  reg [31:0] _RAND_1183;
  reg [31:0] _RAND_1184;
  reg [31:0] _RAND_1185;
  reg [31:0] _RAND_1186;
  reg [31:0] _RAND_1187;
  reg [31:0] _RAND_1188;
  reg [31:0] _RAND_1189;
  reg [31:0] _RAND_1190;
  reg [31:0] _RAND_1191;
  reg [31:0] _RAND_1192;
  reg [31:0] _RAND_1193;
  reg [31:0] _RAND_1194;
  reg [31:0] _RAND_1195;
  reg [31:0] _RAND_1196;
  reg [31:0] _RAND_1197;
  reg [31:0] _RAND_1198;
  reg [31:0] _RAND_1199;
  reg [31:0] _RAND_1200;
  reg [31:0] _RAND_1201;
  reg [31:0] _RAND_1202;
  reg [31:0] _RAND_1203;
  reg [31:0] _RAND_1204;
  reg [31:0] _RAND_1205;
  reg [31:0] _RAND_1206;
  reg [31:0] _RAND_1207;
  reg [31:0] _RAND_1208;
  reg [31:0] _RAND_1209;
  reg [31:0] _RAND_1210;
  reg [31:0] _RAND_1211;
  reg [31:0] _RAND_1212;
  reg [31:0] _RAND_1213;
  reg [31:0] _RAND_1214;
  reg [31:0] _RAND_1215;
  reg [31:0] _RAND_1216;
  reg [31:0] _RAND_1217;
  reg [31:0] _RAND_1218;
  reg [31:0] _RAND_1219;
  reg [31:0] _RAND_1220;
  reg [31:0] _RAND_1221;
  reg [31:0] _RAND_1222;
  reg [31:0] _RAND_1223;
  reg [31:0] _RAND_1224;
  reg [31:0] _RAND_1225;
  reg [31:0] _RAND_1226;
  reg [31:0] _RAND_1227;
  reg [31:0] _RAND_1228;
  reg [31:0] _RAND_1229;
  reg [31:0] _RAND_1230;
  reg [31:0] _RAND_1231;
  reg [31:0] _RAND_1232;
  reg [31:0] _RAND_1233;
  reg [31:0] _RAND_1234;
  reg [31:0] _RAND_1235;
  reg [31:0] _RAND_1236;
  reg [31:0] _RAND_1237;
  reg [31:0] _RAND_1238;
  reg [31:0] _RAND_1239;
  reg [31:0] _RAND_1240;
  reg [31:0] _RAND_1241;
  reg [31:0] _RAND_1242;
  reg [31:0] _RAND_1243;
  reg [31:0] _RAND_1244;
  reg [31:0] _RAND_1245;
  reg [31:0] _RAND_1246;
  reg [31:0] _RAND_1247;
  reg [31:0] _RAND_1248;
  reg [31:0] _RAND_1249;
  reg [31:0] _RAND_1250;
  reg [31:0] _RAND_1251;
  reg [31:0] _RAND_1252;
  reg [31:0] _RAND_1253;
  reg [31:0] _RAND_1254;
  reg [31:0] _RAND_1255;
  reg [31:0] _RAND_1256;
  reg [31:0] _RAND_1257;
  reg [31:0] _RAND_1258;
  reg [31:0] _RAND_1259;
  reg [31:0] _RAND_1260;
  reg [31:0] _RAND_1261;
  reg [31:0] _RAND_1262;
  reg [31:0] _RAND_1263;
  reg [31:0] _RAND_1264;
  reg [31:0] _RAND_1265;
  reg [31:0] _RAND_1266;
  reg [31:0] _RAND_1267;
  reg [31:0] _RAND_1268;
  reg [31:0] _RAND_1269;
  reg [31:0] _RAND_1270;
  reg [31:0] _RAND_1271;
  reg [31:0] _RAND_1272;
  reg [31:0] _RAND_1273;
  reg [31:0] _RAND_1274;
  reg [31:0] _RAND_1275;
  reg [31:0] _RAND_1276;
  reg [31:0] _RAND_1277;
  reg [31:0] _RAND_1278;
  reg [31:0] _RAND_1279;
  reg [31:0] _RAND_1280;
  reg [31:0] _RAND_1281;
  reg [31:0] _RAND_1282;
  reg [31:0] _RAND_1283;
  reg [31:0] _RAND_1284;
  reg [31:0] _RAND_1285;
  reg [31:0] _RAND_1286;
  reg [31:0] _RAND_1287;
  reg [31:0] _RAND_1288;
  reg [31:0] _RAND_1289;
  reg [31:0] _RAND_1290;
  reg [31:0] _RAND_1291;
  reg [31:0] _RAND_1292;
  reg [31:0] _RAND_1293;
  reg [31:0] _RAND_1294;
  reg [31:0] _RAND_1295;
  reg [31:0] _RAND_1296;
  reg [31:0] _RAND_1297;
  reg [31:0] _RAND_1298;
  reg [31:0] _RAND_1299;
  reg [31:0] _RAND_1300;
  reg [31:0] _RAND_1301;
  reg [31:0] _RAND_1302;
  reg [31:0] _RAND_1303;
  reg [31:0] _RAND_1304;
  reg [31:0] _RAND_1305;
  reg [31:0] _RAND_1306;
  reg [31:0] _RAND_1307;
  reg [31:0] _RAND_1308;
  reg [31:0] _RAND_1309;
  reg [31:0] _RAND_1310;
  reg [31:0] _RAND_1311;
  reg [31:0] _RAND_1312;
  reg [31:0] _RAND_1313;
  reg [31:0] _RAND_1314;
  reg [31:0] _RAND_1315;
  reg [31:0] _RAND_1316;
  reg [31:0] _RAND_1317;
  reg [31:0] _RAND_1318;
  reg [31:0] _RAND_1319;
  reg [31:0] _RAND_1320;
  reg [31:0] _RAND_1321;
  reg [31:0] _RAND_1322;
  reg [31:0] _RAND_1323;
  reg [31:0] _RAND_1324;
  reg [31:0] _RAND_1325;
  reg [31:0] _RAND_1326;
  reg [31:0] _RAND_1327;
  reg [31:0] _RAND_1328;
  reg [31:0] _RAND_1329;
  reg [31:0] _RAND_1330;
  reg [31:0] _RAND_1331;
  reg [31:0] _RAND_1332;
  reg [31:0] _RAND_1333;
  reg [31:0] _RAND_1334;
  reg [31:0] _RAND_1335;
  reg [31:0] _RAND_1336;
  reg [31:0] _RAND_1337;
  reg [31:0] _RAND_1338;
  reg [31:0] _RAND_1339;
  reg [31:0] _RAND_1340;
  reg [31:0] _RAND_1341;
  reg [31:0] _RAND_1342;
  reg [31:0] _RAND_1343;
  reg [31:0] _RAND_1344;
  reg [31:0] _RAND_1345;
  reg [31:0] _RAND_1346;
  reg [31:0] _RAND_1347;
  reg [31:0] _RAND_1348;
  reg [31:0] _RAND_1349;
  reg [31:0] _RAND_1350;
  reg [31:0] _RAND_1351;
  reg [31:0] _RAND_1352;
  reg [31:0] _RAND_1353;
  reg [31:0] _RAND_1354;
  reg [31:0] _RAND_1355;
  reg [31:0] _RAND_1356;
  reg [31:0] _RAND_1357;
  reg [31:0] _RAND_1358;
  reg [31:0] _RAND_1359;
  reg [31:0] _RAND_1360;
  reg [31:0] _RAND_1361;
  reg [31:0] _RAND_1362;
  reg [31:0] _RAND_1363;
  reg [31:0] _RAND_1364;
  reg [31:0] _RAND_1365;
  reg [31:0] _RAND_1366;
  reg [31:0] _RAND_1367;
  reg [31:0] _RAND_1368;
  reg [31:0] _RAND_1369;
  reg [31:0] _RAND_1370;
  reg [31:0] _RAND_1371;
  reg [31:0] _RAND_1372;
  reg [31:0] _RAND_1373;
  reg [31:0] _RAND_1374;
  reg [31:0] _RAND_1375;
  reg [31:0] _RAND_1376;
  reg [31:0] _RAND_1377;
  reg [31:0] _RAND_1378;
  reg [31:0] _RAND_1379;
  reg [31:0] _RAND_1380;
  reg [31:0] _RAND_1381;
  reg [31:0] _RAND_1382;
  reg [31:0] _RAND_1383;
  reg [31:0] _RAND_1384;
  reg [31:0] _RAND_1385;
  reg [31:0] _RAND_1386;
  reg [31:0] _RAND_1387;
  reg [31:0] _RAND_1388;
  reg [31:0] _RAND_1389;
  reg [31:0] _RAND_1390;
  reg [31:0] _RAND_1391;
  reg [31:0] _RAND_1392;
  reg [31:0] _RAND_1393;
  reg [31:0] _RAND_1394;
  reg [31:0] _RAND_1395;
  reg [31:0] _RAND_1396;
  reg [31:0] _RAND_1397;
  reg [31:0] _RAND_1398;
  reg [31:0] _RAND_1399;
  reg [31:0] _RAND_1400;
  reg [31:0] _RAND_1401;
  reg [31:0] _RAND_1402;
  reg [31:0] _RAND_1403;
  reg [31:0] _RAND_1404;
  reg [31:0] _RAND_1405;
  reg [31:0] _RAND_1406;
  reg [31:0] _RAND_1407;
  reg [31:0] _RAND_1408;
  reg [31:0] _RAND_1409;
  reg [31:0] _RAND_1410;
  reg [31:0] _RAND_1411;
  reg [31:0] _RAND_1412;
  reg [31:0] _RAND_1413;
  reg [31:0] _RAND_1414;
  reg [31:0] _RAND_1415;
  reg [31:0] _RAND_1416;
  reg [31:0] _RAND_1417;
  reg [31:0] _RAND_1418;
  reg [31:0] _RAND_1419;
  reg [31:0] _RAND_1420;
  reg [31:0] _RAND_1421;
  reg [31:0] _RAND_1422;
  reg [31:0] _RAND_1423;
  reg [31:0] _RAND_1424;
  reg [31:0] _RAND_1425;
  reg [31:0] _RAND_1426;
  reg [31:0] _RAND_1427;
  reg [31:0] _RAND_1428;
  reg [31:0] _RAND_1429;
  reg [31:0] _RAND_1430;
  reg [31:0] _RAND_1431;
  reg [31:0] _RAND_1432;
  reg [31:0] _RAND_1433;
  reg [31:0] _RAND_1434;
  reg [31:0] _RAND_1435;
  reg [31:0] _RAND_1436;
  reg [31:0] _RAND_1437;
  reg [31:0] _RAND_1438;
  reg [31:0] _RAND_1439;
  reg [31:0] _RAND_1440;
  reg [31:0] _RAND_1441;
  reg [31:0] _RAND_1442;
  reg [31:0] _RAND_1443;
  reg [31:0] _RAND_1444;
  reg [31:0] _RAND_1445;
  reg [31:0] _RAND_1446;
  reg [31:0] _RAND_1447;
  reg [31:0] _RAND_1448;
  reg [31:0] _RAND_1449;
  reg [31:0] _RAND_1450;
  reg [31:0] _RAND_1451;
  reg [31:0] _RAND_1452;
  reg [31:0] _RAND_1453;
  reg [31:0] _RAND_1454;
  reg [31:0] _RAND_1455;
  reg [31:0] _RAND_1456;
  reg [31:0] _RAND_1457;
  reg [31:0] _RAND_1458;
  reg [31:0] _RAND_1459;
  reg [31:0] _RAND_1460;
  reg [31:0] _RAND_1461;
  reg [31:0] _RAND_1462;
  reg [31:0] _RAND_1463;
  reg [31:0] _RAND_1464;
  reg [31:0] _RAND_1465;
  reg [31:0] _RAND_1466;
  reg [31:0] _RAND_1467;
  reg [31:0] _RAND_1468;
  reg [31:0] _RAND_1469;
  reg [31:0] _RAND_1470;
  reg [31:0] _RAND_1471;
  reg [31:0] _RAND_1472;
  reg [31:0] _RAND_1473;
  reg [31:0] _RAND_1474;
  reg [31:0] _RAND_1475;
  reg [31:0] _RAND_1476;
  reg [31:0] _RAND_1477;
  reg [31:0] _RAND_1478;
  reg [31:0] _RAND_1479;
  reg [31:0] _RAND_1480;
  reg [31:0] _RAND_1481;
  reg [31:0] _RAND_1482;
  reg [31:0] _RAND_1483;
  reg [31:0] _RAND_1484;
  reg [31:0] _RAND_1485;
  reg [31:0] _RAND_1486;
  reg [31:0] _RAND_1487;
  reg [31:0] _RAND_1488;
  reg [31:0] _RAND_1489;
  reg [31:0] _RAND_1490;
  reg [31:0] _RAND_1491;
  reg [31:0] _RAND_1492;
  reg [31:0] _RAND_1493;
  reg [31:0] _RAND_1494;
  reg [31:0] _RAND_1495;
  reg [31:0] _RAND_1496;
  reg [31:0] _RAND_1497;
  reg [31:0] _RAND_1498;
  reg [31:0] _RAND_1499;
  reg [31:0] _RAND_1500;
  reg [31:0] _RAND_1501;
  reg [31:0] _RAND_1502;
  reg [31:0] _RAND_1503;
  reg [31:0] _RAND_1504;
  reg [31:0] _RAND_1505;
  reg [31:0] _RAND_1506;
  reg [31:0] _RAND_1507;
  reg [31:0] _RAND_1508;
  reg [31:0] _RAND_1509;
  reg [31:0] _RAND_1510;
  reg [31:0] _RAND_1511;
  reg [31:0] _RAND_1512;
  reg [31:0] _RAND_1513;
  reg [31:0] _RAND_1514;
  reg [31:0] _RAND_1515;
  reg [31:0] _RAND_1516;
  reg [31:0] _RAND_1517;
  reg [31:0] _RAND_1518;
  reg [31:0] _RAND_1519;
  reg [31:0] _RAND_1520;
  reg [31:0] _RAND_1521;
  reg [31:0] _RAND_1522;
  reg [31:0] _RAND_1523;
  reg [31:0] _RAND_1524;
  reg [31:0] _RAND_1525;
  reg [31:0] _RAND_1526;
  reg [31:0] _RAND_1527;
  reg [31:0] _RAND_1528;
  reg [31:0] _RAND_1529;
  reg [31:0] _RAND_1530;
  reg [31:0] _RAND_1531;
  reg [31:0] _RAND_1532;
  reg [31:0] _RAND_1533;
  reg [31:0] _RAND_1534;
  reg [31:0] _RAND_1535;
  reg [31:0] _RAND_1536;
  reg [31:0] _RAND_1537;
  reg [31:0] _RAND_1538;
  reg [31:0] _RAND_1539;
  reg [31:0] _RAND_1540;
  reg [31:0] _RAND_1541;
  reg [31:0] _RAND_1542;
  reg [31:0] _RAND_1543;
  reg [31:0] _RAND_1544;
  reg [31:0] _RAND_1545;
  reg [31:0] _RAND_1546;
  reg [31:0] _RAND_1547;
  reg [31:0] _RAND_1548;
  reg [31:0] _RAND_1549;
  reg [31:0] _RAND_1550;
  reg [31:0] _RAND_1551;
  reg [31:0] _RAND_1552;
  reg [31:0] _RAND_1553;
  reg [31:0] _RAND_1554;
  reg [31:0] _RAND_1555;
  reg [31:0] _RAND_1556;
  reg [31:0] _RAND_1557;
  reg [31:0] _RAND_1558;
  reg [31:0] _RAND_1559;
  reg [31:0] _RAND_1560;
  reg [31:0] _RAND_1561;
  reg [31:0] _RAND_1562;
  reg [31:0] _RAND_1563;
  reg [31:0] _RAND_1564;
  reg [31:0] _RAND_1565;
  reg [31:0] _RAND_1566;
  reg [31:0] _RAND_1567;
  reg [31:0] _RAND_1568;
  reg [31:0] _RAND_1569;
  reg [31:0] _RAND_1570;
  reg [31:0] _RAND_1571;
  reg [31:0] _RAND_1572;
  reg [31:0] _RAND_1573;
  reg [31:0] _RAND_1574;
  reg [31:0] _RAND_1575;
  reg [31:0] _RAND_1576;
  reg [31:0] _RAND_1577;
  reg [31:0] _RAND_1578;
  reg [31:0] _RAND_1579;
  reg [31:0] _RAND_1580;
  reg [31:0] _RAND_1581;
  reg [31:0] _RAND_1582;
  reg [31:0] _RAND_1583;
  reg [31:0] _RAND_1584;
  reg [31:0] _RAND_1585;
  reg [31:0] _RAND_1586;
  reg [31:0] _RAND_1587;
  reg [31:0] _RAND_1588;
  reg [31:0] _RAND_1589;
  reg [31:0] _RAND_1590;
  reg [31:0] _RAND_1591;
  reg [31:0] _RAND_1592;
  reg [31:0] _RAND_1593;
  reg [31:0] _RAND_1594;
  reg [31:0] _RAND_1595;
  reg [31:0] _RAND_1596;
  reg [31:0] _RAND_1597;
  reg [31:0] _RAND_1598;
  reg [31:0] _RAND_1599;
  reg [31:0] _RAND_1600;
  reg [31:0] _RAND_1601;
  reg [31:0] _RAND_1602;
  reg [31:0] _RAND_1603;
  reg [31:0] _RAND_1604;
  reg [31:0] _RAND_1605;
  reg [31:0] _RAND_1606;
  reg [31:0] _RAND_1607;
  reg [31:0] _RAND_1608;
  reg [31:0] _RAND_1609;
  reg [31:0] _RAND_1610;
  reg [31:0] _RAND_1611;
  reg [31:0] _RAND_1612;
  reg [31:0] _RAND_1613;
  reg [31:0] _RAND_1614;
  reg [31:0] _RAND_1615;
  reg [31:0] _RAND_1616;
  reg [31:0] _RAND_1617;
  reg [31:0] _RAND_1618;
  reg [31:0] _RAND_1619;
  reg [31:0] _RAND_1620;
  reg [31:0] _RAND_1621;
  reg [31:0] _RAND_1622;
  reg [31:0] _RAND_1623;
  reg [31:0] _RAND_1624;
  reg [31:0] _RAND_1625;
  reg [31:0] _RAND_1626;
  reg [31:0] _RAND_1627;
  reg [31:0] _RAND_1628;
  reg [31:0] _RAND_1629;
  reg [31:0] _RAND_1630;
  reg [31:0] _RAND_1631;
  reg [31:0] _RAND_1632;
  reg [31:0] _RAND_1633;
  reg [31:0] _RAND_1634;
  reg [31:0] _RAND_1635;
  reg [31:0] _RAND_1636;
  reg [31:0] _RAND_1637;
  reg [31:0] _RAND_1638;
  reg [31:0] _RAND_1639;
  reg [31:0] _RAND_1640;
  reg [31:0] _RAND_1641;
  reg [31:0] _RAND_1642;
  reg [31:0] _RAND_1643;
  reg [31:0] _RAND_1644;
  reg [31:0] _RAND_1645;
  reg [31:0] _RAND_1646;
  reg [31:0] _RAND_1647;
  reg [31:0] _RAND_1648;
  reg [31:0] _RAND_1649;
  reg [31:0] _RAND_1650;
  reg [31:0] _RAND_1651;
  reg [31:0] _RAND_1652;
  reg [31:0] _RAND_1653;
  reg [31:0] _RAND_1654;
  reg [31:0] _RAND_1655;
  reg [31:0] _RAND_1656;
  reg [31:0] _RAND_1657;
  reg [31:0] _RAND_1658;
  reg [31:0] _RAND_1659;
  reg [31:0] _RAND_1660;
  reg [31:0] _RAND_1661;
  reg [31:0] _RAND_1662;
  reg [31:0] _RAND_1663;
  reg [31:0] _RAND_1664;
  reg [31:0] _RAND_1665;
  reg [31:0] _RAND_1666;
  reg [31:0] _RAND_1667;
  reg [31:0] _RAND_1668;
  reg [31:0] _RAND_1669;
  reg [31:0] _RAND_1670;
  reg [31:0] _RAND_1671;
  reg [31:0] _RAND_1672;
  reg [31:0] _RAND_1673;
  reg [31:0] _RAND_1674;
  reg [31:0] _RAND_1675;
  reg [31:0] _RAND_1676;
  reg [31:0] _RAND_1677;
  reg [31:0] _RAND_1678;
  reg [31:0] _RAND_1679;
  reg [31:0] _RAND_1680;
  reg [31:0] _RAND_1681;
  reg [31:0] _RAND_1682;
  reg [31:0] _RAND_1683;
  reg [31:0] _RAND_1684;
  reg [31:0] _RAND_1685;
  reg [31:0] _RAND_1686;
  reg [31:0] _RAND_1687;
  reg [31:0] _RAND_1688;
  reg [31:0] _RAND_1689;
  reg [31:0] _RAND_1690;
  reg [31:0] _RAND_1691;
  reg [31:0] _RAND_1692;
  reg [31:0] _RAND_1693;
  reg [31:0] _RAND_1694;
  reg [31:0] _RAND_1695;
  reg [31:0] _RAND_1696;
  reg [31:0] _RAND_1697;
  reg [31:0] _RAND_1698;
  reg [31:0] _RAND_1699;
  reg [31:0] _RAND_1700;
  reg [31:0] _RAND_1701;
  reg [31:0] _RAND_1702;
  reg [31:0] _RAND_1703;
  reg [31:0] _RAND_1704;
  reg [31:0] _RAND_1705;
  reg [31:0] _RAND_1706;
  reg [31:0] _RAND_1707;
  reg [31:0] _RAND_1708;
  reg [31:0] _RAND_1709;
  reg [31:0] _RAND_1710;
  reg [31:0] _RAND_1711;
  reg [31:0] _RAND_1712;
  reg [31:0] _RAND_1713;
  reg [31:0] _RAND_1714;
  reg [31:0] _RAND_1715;
  reg [31:0] _RAND_1716;
  reg [31:0] _RAND_1717;
  reg [31:0] _RAND_1718;
  reg [31:0] _RAND_1719;
  reg [31:0] _RAND_1720;
  reg [31:0] _RAND_1721;
  reg [31:0] _RAND_1722;
  reg [31:0] _RAND_1723;
  reg [31:0] _RAND_1724;
  reg [31:0] _RAND_1725;
  reg [31:0] _RAND_1726;
  reg [31:0] _RAND_1727;
  reg [31:0] _RAND_1728;
  reg [31:0] _RAND_1729;
  reg [31:0] _RAND_1730;
  reg [31:0] _RAND_1731;
  reg [31:0] _RAND_1732;
  reg [31:0] _RAND_1733;
  reg [31:0] _RAND_1734;
  reg [31:0] _RAND_1735;
  reg [31:0] _RAND_1736;
  reg [31:0] _RAND_1737;
  reg [31:0] _RAND_1738;
  reg [31:0] _RAND_1739;
  reg [31:0] _RAND_1740;
  reg [31:0] _RAND_1741;
  reg [31:0] _RAND_1742;
  reg [31:0] _RAND_1743;
  reg [31:0] _RAND_1744;
  reg [31:0] _RAND_1745;
  reg [31:0] _RAND_1746;
  reg [31:0] _RAND_1747;
  reg [31:0] _RAND_1748;
  reg [31:0] _RAND_1749;
  reg [31:0] _RAND_1750;
  reg [31:0] _RAND_1751;
  reg [31:0] _RAND_1752;
  reg [31:0] _RAND_1753;
  reg [31:0] _RAND_1754;
  reg [31:0] _RAND_1755;
  reg [31:0] _RAND_1756;
  reg [31:0] _RAND_1757;
  reg [31:0] _RAND_1758;
  reg [31:0] _RAND_1759;
  reg [31:0] _RAND_1760;
  reg [31:0] _RAND_1761;
  reg [31:0] _RAND_1762;
  reg [31:0] _RAND_1763;
  reg [31:0] _RAND_1764;
  reg [31:0] _RAND_1765;
  reg [31:0] _RAND_1766;
  reg [31:0] _RAND_1767;
  reg [31:0] _RAND_1768;
  reg [31:0] _RAND_1769;
  reg [31:0] _RAND_1770;
  reg [31:0] _RAND_1771;
  reg [31:0] _RAND_1772;
  reg [31:0] _RAND_1773;
  reg [31:0] _RAND_1774;
  reg [31:0] _RAND_1775;
  reg [31:0] _RAND_1776;
  reg [31:0] _RAND_1777;
  reg [31:0] _RAND_1778;
  reg [31:0] _RAND_1779;
  reg [31:0] _RAND_1780;
  reg [31:0] _RAND_1781;
  reg [31:0] _RAND_1782;
  reg [31:0] _RAND_1783;
  reg [31:0] _RAND_1784;
  reg [31:0] _RAND_1785;
  reg [31:0] _RAND_1786;
  reg [31:0] _RAND_1787;
  reg [31:0] _RAND_1788;
  reg [31:0] _RAND_1789;
  reg [31:0] _RAND_1790;
  reg [31:0] _RAND_1791;
  reg [31:0] _RAND_1792;
  reg [31:0] _RAND_1793;
  reg [31:0] _RAND_1794;
  reg [31:0] _RAND_1795;
  reg [31:0] _RAND_1796;
  reg [31:0] _RAND_1797;
  reg [31:0] _RAND_1798;
  reg [31:0] _RAND_1799;
  reg [31:0] _RAND_1800;
  reg [31:0] _RAND_1801;
  reg [31:0] _RAND_1802;
  reg [31:0] _RAND_1803;
  reg [31:0] _RAND_1804;
  reg [31:0] _RAND_1805;
  reg [31:0] _RAND_1806;
  reg [31:0] _RAND_1807;
  reg [31:0] _RAND_1808;
  reg [31:0] _RAND_1809;
  reg [31:0] _RAND_1810;
  reg [31:0] _RAND_1811;
  reg [31:0] _RAND_1812;
  reg [31:0] _RAND_1813;
  reg [31:0] _RAND_1814;
  reg [31:0] _RAND_1815;
  reg [31:0] _RAND_1816;
  reg [31:0] _RAND_1817;
  reg [31:0] _RAND_1818;
  reg [31:0] _RAND_1819;
  reg [31:0] _RAND_1820;
  reg [31:0] _RAND_1821;
  reg [31:0] _RAND_1822;
  reg [31:0] _RAND_1823;
  reg [31:0] _RAND_1824;
  reg [31:0] _RAND_1825;
  reg [31:0] _RAND_1826;
  reg [31:0] _RAND_1827;
  reg [31:0] _RAND_1828;
  reg [31:0] _RAND_1829;
  reg [31:0] _RAND_1830;
  reg [31:0] _RAND_1831;
  reg [31:0] _RAND_1832;
  reg [31:0] _RAND_1833;
  reg [31:0] _RAND_1834;
  reg [31:0] _RAND_1835;
  reg [31:0] _RAND_1836;
  reg [31:0] _RAND_1837;
  reg [31:0] _RAND_1838;
  reg [31:0] _RAND_1839;
  reg [31:0] _RAND_1840;
  reg [31:0] _RAND_1841;
  reg [31:0] _RAND_1842;
  reg [31:0] _RAND_1843;
  reg [31:0] _RAND_1844;
  reg [31:0] _RAND_1845;
  reg [31:0] _RAND_1846;
  reg [31:0] _RAND_1847;
  reg [31:0] _RAND_1848;
  reg [31:0] _RAND_1849;
  reg [31:0] _RAND_1850;
  reg [31:0] _RAND_1851;
  reg [31:0] _RAND_1852;
  reg [31:0] _RAND_1853;
  reg [31:0] _RAND_1854;
  reg [31:0] _RAND_1855;
  reg [31:0] _RAND_1856;
  reg [31:0] _RAND_1857;
  reg [31:0] _RAND_1858;
  reg [31:0] _RAND_1859;
  reg [31:0] _RAND_1860;
  reg [31:0] _RAND_1861;
  reg [31:0] _RAND_1862;
  reg [31:0] _RAND_1863;
  reg [31:0] _RAND_1864;
  reg [31:0] _RAND_1865;
  reg [31:0] _RAND_1866;
  reg [31:0] _RAND_1867;
  reg [31:0] _RAND_1868;
  reg [31:0] _RAND_1869;
  reg [31:0] _RAND_1870;
  reg [31:0] _RAND_1871;
  reg [31:0] _RAND_1872;
  reg [31:0] _RAND_1873;
  reg [31:0] _RAND_1874;
  reg [31:0] _RAND_1875;
  reg [31:0] _RAND_1876;
  reg [31:0] _RAND_1877;
  reg [31:0] _RAND_1878;
  reg [31:0] _RAND_1879;
  reg [31:0] _RAND_1880;
  reg [31:0] _RAND_1881;
  reg [31:0] _RAND_1882;
  reg [31:0] _RAND_1883;
  reg [31:0] _RAND_1884;
  reg [31:0] _RAND_1885;
  reg [31:0] _RAND_1886;
  reg [31:0] _RAND_1887;
  reg [31:0] _RAND_1888;
  reg [31:0] _RAND_1889;
  reg [31:0] _RAND_1890;
  reg [31:0] _RAND_1891;
  reg [31:0] _RAND_1892;
  reg [31:0] _RAND_1893;
  reg [31:0] _RAND_1894;
  reg [31:0] _RAND_1895;
  reg [31:0] _RAND_1896;
  reg [31:0] _RAND_1897;
  reg [31:0] _RAND_1898;
  reg [31:0] _RAND_1899;
  reg [31:0] _RAND_1900;
  reg [31:0] _RAND_1901;
  reg [31:0] _RAND_1902;
  reg [31:0] _RAND_1903;
  reg [31:0] _RAND_1904;
  reg [31:0] _RAND_1905;
  reg [31:0] _RAND_1906;
  reg [31:0] _RAND_1907;
  reg [31:0] _RAND_1908;
  reg [31:0] _RAND_1909;
  reg [31:0] _RAND_1910;
  reg [31:0] _RAND_1911;
  reg [31:0] _RAND_1912;
  reg [31:0] _RAND_1913;
  reg [31:0] _RAND_1914;
  reg [31:0] _RAND_1915;
  reg [31:0] _RAND_1916;
  reg [31:0] _RAND_1917;
  reg [31:0] _RAND_1918;
  reg [31:0] _RAND_1919;
  reg [31:0] _RAND_1920;
  reg [31:0] _RAND_1921;
  reg [31:0] _RAND_1922;
  reg [31:0] _RAND_1923;
  reg [31:0] _RAND_1924;
  reg [31:0] _RAND_1925;
  reg [31:0] _RAND_1926;
  reg [31:0] _RAND_1927;
  reg [31:0] _RAND_1928;
  reg [31:0] _RAND_1929;
  reg [31:0] _RAND_1930;
  reg [31:0] _RAND_1931;
  reg [31:0] _RAND_1932;
  reg [31:0] _RAND_1933;
  reg [31:0] _RAND_1934;
  reg [31:0] _RAND_1935;
  reg [31:0] _RAND_1936;
  reg [31:0] _RAND_1937;
  reg [31:0] _RAND_1938;
  reg [31:0] _RAND_1939;
  reg [31:0] _RAND_1940;
  reg [31:0] _RAND_1941;
  reg [31:0] _RAND_1942;
  reg [31:0] _RAND_1943;
  reg [31:0] _RAND_1944;
  reg [31:0] _RAND_1945;
  reg [31:0] _RAND_1946;
  reg [31:0] _RAND_1947;
  reg [31:0] _RAND_1948;
  reg [31:0] _RAND_1949;
  reg [31:0] _RAND_1950;
  reg [31:0] _RAND_1951;
  reg [31:0] _RAND_1952;
  reg [31:0] _RAND_1953;
  reg [31:0] _RAND_1954;
  reg [31:0] _RAND_1955;
  reg [31:0] _RAND_1956;
  reg [31:0] _RAND_1957;
  reg [31:0] _RAND_1958;
  reg [31:0] _RAND_1959;
  reg [31:0] _RAND_1960;
  reg [31:0] _RAND_1961;
  reg [31:0] _RAND_1962;
  reg [31:0] _RAND_1963;
  reg [31:0] _RAND_1964;
  reg [31:0] _RAND_1965;
  reg [31:0] _RAND_1966;
  reg [31:0] _RAND_1967;
  reg [31:0] _RAND_1968;
  reg [31:0] _RAND_1969;
  reg [31:0] _RAND_1970;
  reg [31:0] _RAND_1971;
  reg [31:0] _RAND_1972;
  reg [31:0] _RAND_1973;
  reg [31:0] _RAND_1974;
  reg [31:0] _RAND_1975;
  reg [31:0] _RAND_1976;
  reg [31:0] _RAND_1977;
  reg [31:0] _RAND_1978;
  reg [31:0] _RAND_1979;
  reg [31:0] _RAND_1980;
  reg [31:0] _RAND_1981;
  reg [31:0] _RAND_1982;
  reg [31:0] _RAND_1983;
  reg [31:0] _RAND_1984;
  reg [31:0] _RAND_1985;
  reg [31:0] _RAND_1986;
  reg [31:0] _RAND_1987;
  reg [31:0] _RAND_1988;
  reg [31:0] _RAND_1989;
  reg [31:0] _RAND_1990;
  reg [31:0] _RAND_1991;
  reg [31:0] _RAND_1992;
  reg [31:0] _RAND_1993;
  reg [31:0] _RAND_1994;
  reg [31:0] _RAND_1995;
  reg [31:0] _RAND_1996;
  reg [31:0] _RAND_1997;
  reg [31:0] _RAND_1998;
  reg [31:0] _RAND_1999;
  reg [31:0] _RAND_2000;
  reg [31:0] _RAND_2001;
  reg [31:0] _RAND_2002;
  reg [31:0] _RAND_2003;
  reg [31:0] _RAND_2004;
  reg [31:0] _RAND_2005;
  reg [31:0] _RAND_2006;
  reg [31:0] _RAND_2007;
  reg [31:0] _RAND_2008;
  reg [31:0] _RAND_2009;
  reg [31:0] _RAND_2010;
  reg [31:0] _RAND_2011;
  reg [31:0] _RAND_2012;
  reg [31:0] _RAND_2013;
  reg [31:0] _RAND_2014;
  reg [31:0] _RAND_2015;
  reg [31:0] _RAND_2016;
  reg [31:0] _RAND_2017;
  reg [31:0] _RAND_2018;
  reg [31:0] _RAND_2019;
  reg [31:0] _RAND_2020;
  reg [31:0] _RAND_2021;
  reg [31:0] _RAND_2022;
  reg [31:0] _RAND_2023;
  reg [31:0] _RAND_2024;
  reg [31:0] _RAND_2025;
  reg [31:0] _RAND_2026;
  reg [31:0] _RAND_2027;
  reg [31:0] _RAND_2028;
  reg [31:0] _RAND_2029;
  reg [31:0] _RAND_2030;
  reg [31:0] _RAND_2031;
  reg [31:0] _RAND_2032;
  reg [31:0] _RAND_2033;
  reg [31:0] _RAND_2034;
  reg [31:0] _RAND_2035;
  reg [31:0] _RAND_2036;
  reg [31:0] _RAND_2037;
  reg [31:0] _RAND_2038;
  reg [31:0] _RAND_2039;
  reg [31:0] _RAND_2040;
  reg [31:0] _RAND_2041;
  reg [31:0] _RAND_2042;
  reg [31:0] _RAND_2043;
  reg [31:0] _RAND_2044;
  reg [31:0] _RAND_2045;
  reg [31:0] _RAND_2046;
  reg [31:0] _RAND_2047;
  reg [31:0] _RAND_2048;
  reg [31:0] _RAND_2049;
  reg [31:0] _RAND_2050;
  reg [31:0] _RAND_2051;
  reg [31:0] _RAND_2052;
  reg [31:0] _RAND_2053;
  reg [31:0] _RAND_2054;
  reg [31:0] _RAND_2055;
  reg [31:0] _RAND_2056;
  reg [31:0] _RAND_2057;
  reg [31:0] _RAND_2058;
  reg [31:0] _RAND_2059;
  reg [31:0] _RAND_2060;
  reg [31:0] _RAND_2061;
  reg [31:0] _RAND_2062;
  reg [31:0] _RAND_2063;
  reg [31:0] _RAND_2064;
  reg [31:0] _RAND_2065;
  reg [31:0] _RAND_2066;
  reg [31:0] _RAND_2067;
  reg [31:0] _RAND_2068;
  reg [31:0] _RAND_2069;
  reg [31:0] _RAND_2070;
  reg [31:0] _RAND_2071;
  reg [31:0] _RAND_2072;
  reg [31:0] _RAND_2073;
  reg [31:0] _RAND_2074;
  reg [31:0] _RAND_2075;
  reg [31:0] _RAND_2076;
  reg [31:0] _RAND_2077;
  reg [31:0] _RAND_2078;
  reg [31:0] _RAND_2079;
  reg [31:0] _RAND_2080;
  reg [31:0] _RAND_2081;
  reg [31:0] _RAND_2082;
  reg [31:0] _RAND_2083;
  reg [31:0] _RAND_2084;
  reg [31:0] _RAND_2085;
  reg [31:0] _RAND_2086;
  reg [31:0] _RAND_2087;
  reg [31:0] _RAND_2088;
  reg [31:0] _RAND_2089;
  reg [31:0] _RAND_2090;
  reg [31:0] _RAND_2091;
  reg [31:0] _RAND_2092;
  reg [31:0] _RAND_2093;
  reg [31:0] _RAND_2094;
  reg [31:0] _RAND_2095;
  reg [31:0] _RAND_2096;
  reg [31:0] _RAND_2097;
  reg [31:0] _RAND_2098;
  reg [31:0] _RAND_2099;
  reg [31:0] _RAND_2100;
  reg [31:0] _RAND_2101;
  reg [31:0] _RAND_2102;
  reg [31:0] _RAND_2103;
  reg [31:0] _RAND_2104;
  reg [31:0] _RAND_2105;
  reg [31:0] _RAND_2106;
  reg [31:0] _RAND_2107;
  reg [31:0] _RAND_2108;
  reg [31:0] _RAND_2109;
  reg [31:0] _RAND_2110;
  reg [31:0] _RAND_2111;
  reg [31:0] _RAND_2112;
  reg [31:0] _RAND_2113;
  reg [31:0] _RAND_2114;
  reg [31:0] _RAND_2115;
  reg [31:0] _RAND_2116;
  reg [31:0] _RAND_2117;
  reg [31:0] _RAND_2118;
  reg [31:0] _RAND_2119;
  reg [31:0] _RAND_2120;
  reg [31:0] _RAND_2121;
  reg [31:0] _RAND_2122;
  reg [31:0] _RAND_2123;
  reg [31:0] _RAND_2124;
  reg [31:0] _RAND_2125;
  reg [31:0] _RAND_2126;
  reg [31:0] _RAND_2127;
  reg [31:0] _RAND_2128;
  reg [31:0] _RAND_2129;
  reg [31:0] _RAND_2130;
  reg [31:0] _RAND_2131;
  reg [31:0] _RAND_2132;
  reg [31:0] _RAND_2133;
  reg [31:0] _RAND_2134;
  reg [31:0] _RAND_2135;
  reg [31:0] _RAND_2136;
  reg [31:0] _RAND_2137;
  reg [31:0] _RAND_2138;
  reg [31:0] _RAND_2139;
  reg [31:0] _RAND_2140;
  reg [31:0] _RAND_2141;
  reg [31:0] _RAND_2142;
  reg [31:0] _RAND_2143;
  reg [31:0] _RAND_2144;
  reg [31:0] _RAND_2145;
  reg [31:0] _RAND_2146;
  reg [31:0] _RAND_2147;
  reg [31:0] _RAND_2148;
  reg [31:0] _RAND_2149;
  reg [31:0] _RAND_2150;
  reg [31:0] _RAND_2151;
  reg [31:0] _RAND_2152;
  reg [31:0] _RAND_2153;
  reg [31:0] _RAND_2154;
  reg [31:0] _RAND_2155;
  reg [31:0] _RAND_2156;
  reg [31:0] _RAND_2157;
  reg [31:0] _RAND_2158;
  reg [31:0] _RAND_2159;
  reg [31:0] _RAND_2160;
  reg [31:0] _RAND_2161;
  reg [31:0] _RAND_2162;
  reg [31:0] _RAND_2163;
  reg [31:0] _RAND_2164;
  reg [31:0] _RAND_2165;
  reg [31:0] _RAND_2166;
  reg [31:0] _RAND_2167;
  reg [31:0] _RAND_2168;
  reg [31:0] _RAND_2169;
  reg [31:0] _RAND_2170;
  reg [31:0] _RAND_2171;
  reg [31:0] _RAND_2172;
  reg [31:0] _RAND_2173;
  reg [31:0] _RAND_2174;
  reg [31:0] _RAND_2175;
  reg [31:0] _RAND_2176;
  reg [31:0] _RAND_2177;
  reg [31:0] _RAND_2178;
  reg [31:0] _RAND_2179;
  reg [31:0] _RAND_2180;
  reg [31:0] _RAND_2181;
  reg [31:0] _RAND_2182;
  reg [31:0] _RAND_2183;
  reg [31:0] _RAND_2184;
  reg [31:0] _RAND_2185;
  reg [31:0] _RAND_2186;
  reg [31:0] _RAND_2187;
  reg [31:0] _RAND_2188;
  reg [31:0] _RAND_2189;
  reg [31:0] _RAND_2190;
  reg [31:0] _RAND_2191;
  reg [31:0] _RAND_2192;
  reg [31:0] _RAND_2193;
  reg [31:0] _RAND_2194;
  reg [31:0] _RAND_2195;
  reg [31:0] _RAND_2196;
  reg [31:0] _RAND_2197;
  reg [31:0] _RAND_2198;
  reg [31:0] _RAND_2199;
  reg [31:0] _RAND_2200;
  reg [31:0] _RAND_2201;
  reg [31:0] _RAND_2202;
  reg [31:0] _RAND_2203;
  reg [31:0] _RAND_2204;
  reg [31:0] _RAND_2205;
  reg [31:0] _RAND_2206;
  reg [31:0] _RAND_2207;
  reg [31:0] _RAND_2208;
  reg [31:0] _RAND_2209;
  reg [31:0] _RAND_2210;
  reg [31:0] _RAND_2211;
  reg [31:0] _RAND_2212;
  reg [31:0] _RAND_2213;
  reg [31:0] _RAND_2214;
  reg [31:0] _RAND_2215;
  reg [31:0] _RAND_2216;
  reg [31:0] _RAND_2217;
  reg [31:0] _RAND_2218;
  reg [31:0] _RAND_2219;
  reg [31:0] _RAND_2220;
  reg [31:0] _RAND_2221;
  reg [31:0] _RAND_2222;
  reg [31:0] _RAND_2223;
  reg [31:0] _RAND_2224;
  reg [31:0] _RAND_2225;
  reg [31:0] _RAND_2226;
  reg [31:0] _RAND_2227;
  reg [31:0] _RAND_2228;
  reg [31:0] _RAND_2229;
  reg [31:0] _RAND_2230;
  reg [31:0] _RAND_2231;
  reg [31:0] _RAND_2232;
  reg [31:0] _RAND_2233;
  reg [31:0] _RAND_2234;
  reg [31:0] _RAND_2235;
  reg [31:0] _RAND_2236;
  reg [31:0] _RAND_2237;
  reg [31:0] _RAND_2238;
  reg [31:0] _RAND_2239;
  reg [31:0] _RAND_2240;
  reg [31:0] _RAND_2241;
  reg [31:0] _RAND_2242;
  reg [31:0] _RAND_2243;
  reg [31:0] _RAND_2244;
  reg [31:0] _RAND_2245;
  reg [31:0] _RAND_2246;
  reg [31:0] _RAND_2247;
  reg [31:0] _RAND_2248;
  reg [31:0] _RAND_2249;
  reg [31:0] _RAND_2250;
  reg [31:0] _RAND_2251;
  reg [31:0] _RAND_2252;
  reg [31:0] _RAND_2253;
  reg [31:0] _RAND_2254;
  reg [31:0] _RAND_2255;
  reg [31:0] _RAND_2256;
  reg [31:0] _RAND_2257;
  reg [31:0] _RAND_2258;
  reg [31:0] _RAND_2259;
  reg [31:0] _RAND_2260;
  reg [31:0] _RAND_2261;
  reg [31:0] _RAND_2262;
  reg [31:0] _RAND_2263;
  reg [31:0] _RAND_2264;
  reg [31:0] _RAND_2265;
  reg [31:0] _RAND_2266;
  reg [31:0] _RAND_2267;
  reg [31:0] _RAND_2268;
  reg [31:0] _RAND_2269;
  reg [31:0] _RAND_2270;
  reg [31:0] _RAND_2271;
  reg [31:0] _RAND_2272;
  reg [31:0] _RAND_2273;
  reg [31:0] _RAND_2274;
  reg [31:0] _RAND_2275;
  reg [31:0] _RAND_2276;
  reg [31:0] _RAND_2277;
  reg [31:0] _RAND_2278;
  reg [31:0] _RAND_2279;
  reg [31:0] _RAND_2280;
  reg [31:0] _RAND_2281;
  reg [31:0] _RAND_2282;
  reg [31:0] _RAND_2283;
  reg [31:0] _RAND_2284;
  reg [31:0] _RAND_2285;
  reg [31:0] _RAND_2286;
  reg [31:0] _RAND_2287;
  reg [31:0] _RAND_2288;
  reg [31:0] _RAND_2289;
  reg [31:0] _RAND_2290;
  reg [31:0] _RAND_2291;
  reg [31:0] _RAND_2292;
  reg [31:0] _RAND_2293;
  reg [31:0] _RAND_2294;
  reg [31:0] _RAND_2295;
  reg [31:0] _RAND_2296;
  reg [31:0] _RAND_2297;
  reg [31:0] _RAND_2298;
  reg [31:0] _RAND_2299;
  reg [31:0] _RAND_2300;
  reg [31:0] _RAND_2301;
  reg [31:0] _RAND_2302;
  reg [31:0] _RAND_2303;
  reg [31:0] _RAND_2304;
  reg [31:0] _RAND_2305;
  reg [31:0] _RAND_2306;
  reg [31:0] _RAND_2307;
  reg [31:0] _RAND_2308;
  reg [31:0] _RAND_2309;
  reg [31:0] _RAND_2310;
  reg [31:0] _RAND_2311;
  reg [31:0] _RAND_2312;
  reg [31:0] _RAND_2313;
  reg [31:0] _RAND_2314;
  reg [31:0] _RAND_2315;
  reg [31:0] _RAND_2316;
  reg [31:0] _RAND_2317;
  reg [31:0] _RAND_2318;
  reg [31:0] _RAND_2319;
  reg [31:0] _RAND_2320;
  reg [31:0] _RAND_2321;
  reg [31:0] _RAND_2322;
  reg [31:0] _RAND_2323;
  reg [31:0] _RAND_2324;
  reg [31:0] _RAND_2325;
  reg [31:0] _RAND_2326;
  reg [31:0] _RAND_2327;
  reg [31:0] _RAND_2328;
  reg [31:0] _RAND_2329;
  reg [31:0] _RAND_2330;
  reg [31:0] _RAND_2331;
  reg [31:0] _RAND_2332;
  reg [31:0] _RAND_2333;
  reg [31:0] _RAND_2334;
  reg [31:0] _RAND_2335;
  reg [31:0] _RAND_2336;
  reg [31:0] _RAND_2337;
  reg [31:0] _RAND_2338;
  reg [31:0] _RAND_2339;
  reg [31:0] _RAND_2340;
  reg [31:0] _RAND_2341;
  reg [31:0] _RAND_2342;
  reg [31:0] _RAND_2343;
  reg [31:0] _RAND_2344;
  reg [31:0] _RAND_2345;
  reg [31:0] _RAND_2346;
  reg [31:0] _RAND_2347;
  reg [31:0] _RAND_2348;
  reg [31:0] _RAND_2349;
  reg [31:0] _RAND_2350;
  reg [31:0] _RAND_2351;
  reg [31:0] _RAND_2352;
  reg [31:0] _RAND_2353;
  reg [31:0] _RAND_2354;
  reg [31:0] _RAND_2355;
  reg [31:0] _RAND_2356;
  reg [31:0] _RAND_2357;
  reg [31:0] _RAND_2358;
  reg [31:0] _RAND_2359;
  reg [31:0] _RAND_2360;
  reg [31:0] _RAND_2361;
  reg [31:0] _RAND_2362;
  reg [31:0] _RAND_2363;
  reg [31:0] _RAND_2364;
  reg [31:0] _RAND_2365;
  reg [31:0] _RAND_2366;
  reg [31:0] _RAND_2367;
  reg [31:0] _RAND_2368;
  reg [31:0] _RAND_2369;
  reg [31:0] _RAND_2370;
  reg [31:0] _RAND_2371;
  reg [31:0] _RAND_2372;
  reg [31:0] _RAND_2373;
  reg [31:0] _RAND_2374;
  reg [31:0] _RAND_2375;
  reg [31:0] _RAND_2376;
  reg [31:0] _RAND_2377;
  reg [31:0] _RAND_2378;
  reg [31:0] _RAND_2379;
  reg [31:0] _RAND_2380;
  reg [31:0] _RAND_2381;
  reg [31:0] _RAND_2382;
  reg [31:0] _RAND_2383;
  reg [31:0] _RAND_2384;
  reg [31:0] _RAND_2385;
  reg [31:0] _RAND_2386;
  reg [31:0] _RAND_2387;
  reg [31:0] _RAND_2388;
  reg [31:0] _RAND_2389;
  reg [31:0] _RAND_2390;
  reg [31:0] _RAND_2391;
  reg [31:0] _RAND_2392;
  reg [31:0] _RAND_2393;
  reg [31:0] _RAND_2394;
  reg [31:0] _RAND_2395;
  reg [31:0] _RAND_2396;
  reg [31:0] _RAND_2397;
  reg [31:0] _RAND_2398;
  reg [31:0] _RAND_2399;
  reg [31:0] _RAND_2400;
  reg [31:0] _RAND_2401;
  reg [31:0] _RAND_2402;
  reg [31:0] _RAND_2403;
  reg [31:0] _RAND_2404;
  reg [31:0] _RAND_2405;
  reg [31:0] _RAND_2406;
  reg [31:0] _RAND_2407;
  reg [31:0] _RAND_2408;
  reg [31:0] _RAND_2409;
  reg [31:0] _RAND_2410;
  reg [31:0] _RAND_2411;
  reg [31:0] _RAND_2412;
  reg [31:0] _RAND_2413;
  reg [31:0] _RAND_2414;
  reg [31:0] _RAND_2415;
  reg [31:0] _RAND_2416;
  reg [31:0] _RAND_2417;
  reg [31:0] _RAND_2418;
  reg [31:0] _RAND_2419;
  reg [31:0] _RAND_2420;
  reg [31:0] _RAND_2421;
  reg [31:0] _RAND_2422;
  reg [31:0] _RAND_2423;
  reg [31:0] _RAND_2424;
  reg [31:0] _RAND_2425;
  reg [31:0] _RAND_2426;
  reg [31:0] _RAND_2427;
  reg [31:0] _RAND_2428;
  reg [31:0] _RAND_2429;
  reg [31:0] _RAND_2430;
  reg [31:0] _RAND_2431;
  reg [31:0] _RAND_2432;
  reg [31:0] _RAND_2433;
  reg [31:0] _RAND_2434;
  reg [31:0] _RAND_2435;
  reg [31:0] _RAND_2436;
  reg [31:0] _RAND_2437;
  reg [31:0] _RAND_2438;
  reg [31:0] _RAND_2439;
  reg [31:0] _RAND_2440;
  reg [31:0] _RAND_2441;
  reg [31:0] _RAND_2442;
  reg [31:0] _RAND_2443;
  reg [31:0] _RAND_2444;
  reg [31:0] _RAND_2445;
  reg [31:0] _RAND_2446;
  reg [31:0] _RAND_2447;
  reg [31:0] _RAND_2448;
  reg [31:0] _RAND_2449;
  reg [31:0] _RAND_2450;
  reg [31:0] _RAND_2451;
  reg [31:0] _RAND_2452;
  reg [31:0] _RAND_2453;
  reg [31:0] _RAND_2454;
  reg [31:0] _RAND_2455;
  reg [31:0] _RAND_2456;
  reg [31:0] _RAND_2457;
  reg [31:0] _RAND_2458;
  reg [31:0] _RAND_2459;
  reg [31:0] _RAND_2460;
  reg [31:0] _RAND_2461;
  reg [31:0] _RAND_2462;
  reg [31:0] _RAND_2463;
  reg [31:0] _RAND_2464;
  reg [31:0] _RAND_2465;
  reg [31:0] _RAND_2466;
  reg [31:0] _RAND_2467;
  reg [31:0] _RAND_2468;
  reg [31:0] _RAND_2469;
  reg [31:0] _RAND_2470;
  reg [31:0] _RAND_2471;
  reg [31:0] _RAND_2472;
  reg [31:0] _RAND_2473;
  reg [31:0] _RAND_2474;
  reg [31:0] _RAND_2475;
  reg [31:0] _RAND_2476;
  reg [31:0] _RAND_2477;
  reg [31:0] _RAND_2478;
  reg [31:0] _RAND_2479;
  reg [31:0] _RAND_2480;
  reg [31:0] _RAND_2481;
  reg [31:0] _RAND_2482;
  reg [31:0] _RAND_2483;
  reg [31:0] _RAND_2484;
  reg [31:0] _RAND_2485;
  reg [31:0] _RAND_2486;
  reg [31:0] _RAND_2487;
  reg [31:0] _RAND_2488;
  reg [31:0] _RAND_2489;
  reg [31:0] _RAND_2490;
  reg [31:0] _RAND_2491;
  reg [31:0] _RAND_2492;
  reg [31:0] _RAND_2493;
  reg [31:0] _RAND_2494;
  reg [31:0] _RAND_2495;
  reg [31:0] _RAND_2496;
  reg [31:0] _RAND_2497;
  reg [31:0] _RAND_2498;
  reg [31:0] _RAND_2499;
  reg [31:0] _RAND_2500;
  reg [31:0] _RAND_2501;
  reg [31:0] _RAND_2502;
  reg [31:0] _RAND_2503;
  reg [31:0] _RAND_2504;
  reg [31:0] _RAND_2505;
  reg [31:0] _RAND_2506;
  reg [31:0] _RAND_2507;
  reg [31:0] _RAND_2508;
  reg [31:0] _RAND_2509;
  reg [31:0] _RAND_2510;
  reg [31:0] _RAND_2511;
  reg [31:0] _RAND_2512;
  reg [31:0] _RAND_2513;
  reg [31:0] _RAND_2514;
  reg [31:0] _RAND_2515;
  reg [31:0] _RAND_2516;
  reg [31:0] _RAND_2517;
  reg [31:0] _RAND_2518;
  reg [31:0] _RAND_2519;
  reg [31:0] _RAND_2520;
  reg [31:0] _RAND_2521;
  reg [31:0] _RAND_2522;
  reg [31:0] _RAND_2523;
  reg [31:0] _RAND_2524;
  reg [31:0] _RAND_2525;
  reg [31:0] _RAND_2526;
  reg [31:0] _RAND_2527;
  reg [31:0] _RAND_2528;
  reg [31:0] _RAND_2529;
  reg [31:0] _RAND_2530;
  reg [31:0] _RAND_2531;
  reg [31:0] _RAND_2532;
  reg [31:0] _RAND_2533;
  reg [31:0] _RAND_2534;
  reg [31:0] _RAND_2535;
  reg [31:0] _RAND_2536;
  reg [31:0] _RAND_2537;
  reg [31:0] _RAND_2538;
  reg [31:0] _RAND_2539;
  reg [31:0] _RAND_2540;
  reg [31:0] _RAND_2541;
  reg [31:0] _RAND_2542;
  reg [31:0] _RAND_2543;
  reg [31:0] _RAND_2544;
  reg [31:0] _RAND_2545;
  reg [31:0] _RAND_2546;
  reg [31:0] _RAND_2547;
  reg [31:0] _RAND_2548;
  reg [31:0] _RAND_2549;
  reg [31:0] _RAND_2550;
  reg [31:0] _RAND_2551;
  reg [31:0] _RAND_2552;
  reg [31:0] _RAND_2553;
  reg [31:0] _RAND_2554;
  reg [31:0] _RAND_2555;
  reg [31:0] _RAND_2556;
  reg [31:0] _RAND_2557;
  reg [31:0] _RAND_2558;
  reg [31:0] _RAND_2559;
  reg [31:0] _RAND_2560;
  reg [31:0] _RAND_2561;
  reg [31:0] _RAND_2562;
  reg [31:0] _RAND_2563;
  reg [31:0] _RAND_2564;
  reg [31:0] _RAND_2565;
  reg [31:0] _RAND_2566;
  reg [31:0] _RAND_2567;
  reg [31:0] _RAND_2568;
  reg [31:0] _RAND_2569;
  reg [31:0] _RAND_2570;
  reg [31:0] _RAND_2571;
  reg [31:0] _RAND_2572;
  reg [31:0] _RAND_2573;
  reg [31:0] _RAND_2574;
  reg [31:0] _RAND_2575;
  reg [31:0] _RAND_2576;
  reg [31:0] _RAND_2577;
  reg [31:0] _RAND_2578;
  reg [31:0] _RAND_2579;
  reg [31:0] _RAND_2580;
  reg [31:0] _RAND_2581;
  reg [31:0] _RAND_2582;
  reg [31:0] _RAND_2583;
  reg [31:0] _RAND_2584;
  reg [31:0] _RAND_2585;
  reg [31:0] _RAND_2586;
  reg [31:0] _RAND_2587;
  reg [31:0] _RAND_2588;
  reg [31:0] _RAND_2589;
  reg [31:0] _RAND_2590;
  reg [31:0] _RAND_2591;
  reg [31:0] _RAND_2592;
  reg [31:0] _RAND_2593;
  reg [31:0] _RAND_2594;
  reg [31:0] _RAND_2595;
  reg [31:0] _RAND_2596;
  reg [31:0] _RAND_2597;
  reg [31:0] _RAND_2598;
  reg [31:0] _RAND_2599;
  reg [31:0] _RAND_2600;
  reg [31:0] _RAND_2601;
  reg [31:0] _RAND_2602;
  reg [31:0] _RAND_2603;
  reg [31:0] _RAND_2604;
  reg [31:0] _RAND_2605;
  reg [31:0] _RAND_2606;
  reg [31:0] _RAND_2607;
  reg [31:0] _RAND_2608;
  reg [31:0] _RAND_2609;
  reg [31:0] _RAND_2610;
  reg [31:0] _RAND_2611;
  reg [31:0] _RAND_2612;
  reg [31:0] _RAND_2613;
  reg [31:0] _RAND_2614;
  reg [31:0] _RAND_2615;
  reg [31:0] _RAND_2616;
  reg [31:0] _RAND_2617;
  reg [31:0] _RAND_2618;
  reg [31:0] _RAND_2619;
  reg [31:0] _RAND_2620;
  reg [31:0] _RAND_2621;
  reg [31:0] _RAND_2622;
  reg [31:0] _RAND_2623;
  reg [31:0] _RAND_2624;
  reg [31:0] _RAND_2625;
  reg [31:0] _RAND_2626;
  reg [31:0] _RAND_2627;
  reg [31:0] _RAND_2628;
  reg [31:0] _RAND_2629;
  reg [31:0] _RAND_2630;
  reg [31:0] _RAND_2631;
  reg [31:0] _RAND_2632;
  reg [31:0] _RAND_2633;
  reg [31:0] _RAND_2634;
  reg [31:0] _RAND_2635;
  reg [31:0] _RAND_2636;
  reg [31:0] _RAND_2637;
  reg [31:0] _RAND_2638;
  reg [31:0] _RAND_2639;
  reg [31:0] _RAND_2640;
  reg [31:0] _RAND_2641;
  reg [31:0] _RAND_2642;
  reg [31:0] _RAND_2643;
  reg [31:0] _RAND_2644;
  reg [31:0] _RAND_2645;
  reg [31:0] _RAND_2646;
  reg [31:0] _RAND_2647;
  reg [31:0] _RAND_2648;
  reg [31:0] _RAND_2649;
  reg [31:0] _RAND_2650;
  reg [31:0] _RAND_2651;
  reg [31:0] _RAND_2652;
  reg [31:0] _RAND_2653;
  reg [31:0] _RAND_2654;
  reg [31:0] _RAND_2655;
  reg [31:0] _RAND_2656;
  reg [31:0] _RAND_2657;
  reg [31:0] _RAND_2658;
  reg [31:0] _RAND_2659;
  reg [31:0] _RAND_2660;
  reg [31:0] _RAND_2661;
  reg [31:0] _RAND_2662;
  reg [31:0] _RAND_2663;
  reg [31:0] _RAND_2664;
  reg [31:0] _RAND_2665;
  reg [31:0] _RAND_2666;
  reg [31:0] _RAND_2667;
  reg [31:0] _RAND_2668;
  reg [31:0] _RAND_2669;
  reg [31:0] _RAND_2670;
  reg [31:0] _RAND_2671;
  reg [31:0] _RAND_2672;
  reg [31:0] _RAND_2673;
  reg [31:0] _RAND_2674;
  reg [31:0] _RAND_2675;
  reg [31:0] _RAND_2676;
  reg [31:0] _RAND_2677;
  reg [31:0] _RAND_2678;
  reg [31:0] _RAND_2679;
  reg [31:0] _RAND_2680;
  reg [31:0] _RAND_2681;
  reg [31:0] _RAND_2682;
  reg [31:0] _RAND_2683;
  reg [31:0] _RAND_2684;
  reg [31:0] _RAND_2685;
  reg [31:0] _RAND_2686;
  reg [31:0] _RAND_2687;
  reg [31:0] _RAND_2688;
  reg [31:0] _RAND_2689;
  reg [31:0] _RAND_2690;
  reg [31:0] _RAND_2691;
  reg [31:0] _RAND_2692;
  reg [31:0] _RAND_2693;
  reg [31:0] _RAND_2694;
  reg [31:0] _RAND_2695;
  reg [31:0] _RAND_2696;
  reg [31:0] _RAND_2697;
  reg [31:0] _RAND_2698;
  reg [31:0] _RAND_2699;
  reg [31:0] _RAND_2700;
  reg [31:0] _RAND_2701;
  reg [31:0] _RAND_2702;
  reg [31:0] _RAND_2703;
  reg [31:0] _RAND_2704;
  reg [31:0] _RAND_2705;
  reg [31:0] _RAND_2706;
  reg [31:0] _RAND_2707;
  reg [31:0] _RAND_2708;
  reg [31:0] _RAND_2709;
  reg [31:0] _RAND_2710;
  reg [31:0] _RAND_2711;
  reg [31:0] _RAND_2712;
  reg [31:0] _RAND_2713;
  reg [31:0] _RAND_2714;
  reg [31:0] _RAND_2715;
  reg [31:0] _RAND_2716;
  reg [31:0] _RAND_2717;
  reg [31:0] _RAND_2718;
  reg [31:0] _RAND_2719;
  reg [31:0] _RAND_2720;
  reg [31:0] _RAND_2721;
  reg [31:0] _RAND_2722;
  reg [31:0] _RAND_2723;
  reg [31:0] _RAND_2724;
  reg [31:0] _RAND_2725;
  reg [31:0] _RAND_2726;
  reg [31:0] _RAND_2727;
  reg [31:0] _RAND_2728;
  reg [31:0] _RAND_2729;
  reg [31:0] _RAND_2730;
  reg [31:0] _RAND_2731;
  reg [31:0] _RAND_2732;
  reg [31:0] _RAND_2733;
  reg [31:0] _RAND_2734;
  reg [31:0] _RAND_2735;
  reg [31:0] _RAND_2736;
  reg [31:0] _RAND_2737;
  reg [31:0] _RAND_2738;
  reg [31:0] _RAND_2739;
  reg [31:0] _RAND_2740;
  reg [31:0] _RAND_2741;
  reg [31:0] _RAND_2742;
  reg [31:0] _RAND_2743;
  reg [31:0] _RAND_2744;
  reg [31:0] _RAND_2745;
  reg [31:0] _RAND_2746;
  reg [31:0] _RAND_2747;
  reg [31:0] _RAND_2748;
  reg [31:0] _RAND_2749;
  reg [31:0] _RAND_2750;
  reg [31:0] _RAND_2751;
  reg [31:0] _RAND_2752;
  reg [31:0] _RAND_2753;
  reg [31:0] _RAND_2754;
  reg [31:0] _RAND_2755;
  reg [31:0] _RAND_2756;
  reg [31:0] _RAND_2757;
  reg [31:0] _RAND_2758;
  reg [31:0] _RAND_2759;
  reg [31:0] _RAND_2760;
  reg [31:0] _RAND_2761;
  reg [31:0] _RAND_2762;
  reg [31:0] _RAND_2763;
  reg [31:0] _RAND_2764;
  reg [31:0] _RAND_2765;
  reg [31:0] _RAND_2766;
  reg [31:0] _RAND_2767;
  reg [31:0] _RAND_2768;
  reg [31:0] _RAND_2769;
  reg [31:0] _RAND_2770;
  reg [31:0] _RAND_2771;
  reg [31:0] _RAND_2772;
  reg [31:0] _RAND_2773;
  reg [31:0] _RAND_2774;
  reg [31:0] _RAND_2775;
  reg [31:0] _RAND_2776;
  reg [31:0] _RAND_2777;
  reg [31:0] _RAND_2778;
  reg [31:0] _RAND_2779;
  reg [31:0] _RAND_2780;
  reg [31:0] _RAND_2781;
  reg [31:0] _RAND_2782;
  reg [31:0] _RAND_2783;
  reg [31:0] _RAND_2784;
  reg [31:0] _RAND_2785;
  reg [31:0] _RAND_2786;
  reg [31:0] _RAND_2787;
  reg [31:0] _RAND_2788;
  reg [31:0] _RAND_2789;
  reg [31:0] _RAND_2790;
  reg [31:0] _RAND_2791;
  reg [31:0] _RAND_2792;
  reg [31:0] _RAND_2793;
  reg [31:0] _RAND_2794;
  reg [31:0] _RAND_2795;
  reg [31:0] _RAND_2796;
  reg [31:0] _RAND_2797;
  reg [31:0] _RAND_2798;
  reg [31:0] _RAND_2799;
  reg [31:0] _RAND_2800;
  reg [31:0] _RAND_2801;
  reg [31:0] _RAND_2802;
  reg [31:0] _RAND_2803;
  reg [31:0] _RAND_2804;
  reg [31:0] _RAND_2805;
  reg [31:0] _RAND_2806;
  reg [31:0] _RAND_2807;
  reg [31:0] _RAND_2808;
  reg [31:0] _RAND_2809;
  reg [31:0] _RAND_2810;
  reg [31:0] _RAND_2811;
  reg [31:0] _RAND_2812;
  reg [31:0] _RAND_2813;
  reg [31:0] _RAND_2814;
  reg [31:0] _RAND_2815;
  reg [31:0] _RAND_2816;
  reg [31:0] _RAND_2817;
  reg [31:0] _RAND_2818;
  reg [31:0] _RAND_2819;
  reg [31:0] _RAND_2820;
  reg [31:0] _RAND_2821;
  reg [31:0] _RAND_2822;
  reg [31:0] _RAND_2823;
  reg [31:0] _RAND_2824;
  reg [31:0] _RAND_2825;
  reg [31:0] _RAND_2826;
  reg [31:0] _RAND_2827;
  reg [31:0] _RAND_2828;
  reg [31:0] _RAND_2829;
  reg [31:0] _RAND_2830;
  reg [31:0] _RAND_2831;
  reg [31:0] _RAND_2832;
  reg [31:0] _RAND_2833;
  reg [31:0] _RAND_2834;
  reg [31:0] _RAND_2835;
  reg [31:0] _RAND_2836;
  reg [31:0] _RAND_2837;
  reg [31:0] _RAND_2838;
  reg [31:0] _RAND_2839;
  reg [31:0] _RAND_2840;
  reg [31:0] _RAND_2841;
  reg [31:0] _RAND_2842;
  reg [31:0] _RAND_2843;
  reg [31:0] _RAND_2844;
  reg [31:0] _RAND_2845;
  reg [31:0] _RAND_2846;
  reg [31:0] _RAND_2847;
  reg [31:0] _RAND_2848;
  reg [31:0] _RAND_2849;
  reg [31:0] _RAND_2850;
  reg [31:0] _RAND_2851;
  reg [31:0] _RAND_2852;
  reg [31:0] _RAND_2853;
  reg [31:0] _RAND_2854;
  reg [31:0] _RAND_2855;
  reg [31:0] _RAND_2856;
  reg [31:0] _RAND_2857;
  reg [31:0] _RAND_2858;
  reg [31:0] _RAND_2859;
  reg [31:0] _RAND_2860;
  reg [31:0] _RAND_2861;
  reg [31:0] _RAND_2862;
  reg [31:0] _RAND_2863;
  reg [31:0] _RAND_2864;
  reg [31:0] _RAND_2865;
  reg [31:0] _RAND_2866;
  reg [31:0] _RAND_2867;
  reg [31:0] _RAND_2868;
  reg [31:0] _RAND_2869;
  reg [31:0] _RAND_2870;
  reg [31:0] _RAND_2871;
  reg [31:0] _RAND_2872;
  reg [31:0] _RAND_2873;
  reg [31:0] _RAND_2874;
  reg [31:0] _RAND_2875;
  reg [31:0] _RAND_2876;
  reg [31:0] _RAND_2877;
  reg [31:0] _RAND_2878;
  reg [31:0] _RAND_2879;
  reg [31:0] _RAND_2880;
  reg [31:0] _RAND_2881;
  reg [31:0] _RAND_2882;
  reg [31:0] _RAND_2883;
  reg [31:0] _RAND_2884;
  reg [31:0] _RAND_2885;
  reg [31:0] _RAND_2886;
  reg [31:0] _RAND_2887;
  reg [31:0] _RAND_2888;
  reg [31:0] _RAND_2889;
  reg [31:0] _RAND_2890;
  reg [31:0] _RAND_2891;
  reg [31:0] _RAND_2892;
  reg [31:0] _RAND_2893;
  reg [31:0] _RAND_2894;
  reg [31:0] _RAND_2895;
  reg [31:0] _RAND_2896;
  reg [31:0] _RAND_2897;
  reg [31:0] _RAND_2898;
  reg [31:0] _RAND_2899;
  reg [31:0] _RAND_2900;
  reg [31:0] _RAND_2901;
  reg [31:0] _RAND_2902;
  reg [31:0] _RAND_2903;
  reg [31:0] _RAND_2904;
  reg [31:0] _RAND_2905;
  reg [31:0] _RAND_2906;
  reg [31:0] _RAND_2907;
  reg [31:0] _RAND_2908;
  reg [31:0] _RAND_2909;
  reg [31:0] _RAND_2910;
  reg [31:0] _RAND_2911;
  reg [31:0] _RAND_2912;
  reg [31:0] _RAND_2913;
  reg [31:0] _RAND_2914;
  reg [31:0] _RAND_2915;
  reg [31:0] _RAND_2916;
  reg [31:0] _RAND_2917;
  reg [31:0] _RAND_2918;
  reg [31:0] _RAND_2919;
  reg [31:0] _RAND_2920;
  reg [31:0] _RAND_2921;
  reg [31:0] _RAND_2922;
  reg [31:0] _RAND_2923;
  reg [31:0] _RAND_2924;
  reg [31:0] _RAND_2925;
  reg [31:0] _RAND_2926;
  reg [31:0] _RAND_2927;
  reg [31:0] _RAND_2928;
  reg [31:0] _RAND_2929;
  reg [31:0] _RAND_2930;
  reg [31:0] _RAND_2931;
  reg [31:0] _RAND_2932;
  reg [31:0] _RAND_2933;
  reg [31:0] _RAND_2934;
  reg [31:0] _RAND_2935;
  reg [31:0] _RAND_2936;
  reg [31:0] _RAND_2937;
  reg [31:0] _RAND_2938;
  reg [31:0] _RAND_2939;
  reg [31:0] _RAND_2940;
  reg [31:0] _RAND_2941;
  reg [31:0] _RAND_2942;
  reg [31:0] _RAND_2943;
  reg [31:0] _RAND_2944;
  reg [31:0] _RAND_2945;
  reg [31:0] _RAND_2946;
  reg [31:0] _RAND_2947;
  reg [31:0] _RAND_2948;
  reg [31:0] _RAND_2949;
  reg [31:0] _RAND_2950;
  reg [31:0] _RAND_2951;
  reg [31:0] _RAND_2952;
  reg [31:0] _RAND_2953;
  reg [31:0] _RAND_2954;
  reg [31:0] _RAND_2955;
  reg [31:0] _RAND_2956;
  reg [31:0] _RAND_2957;
  reg [31:0] _RAND_2958;
  reg [31:0] _RAND_2959;
  reg [31:0] _RAND_2960;
  reg [31:0] _RAND_2961;
  reg [31:0] _RAND_2962;
  reg [31:0] _RAND_2963;
  reg [31:0] _RAND_2964;
  reg [31:0] _RAND_2965;
  reg [31:0] _RAND_2966;
  reg [31:0] _RAND_2967;
  reg [31:0] _RAND_2968;
  reg [31:0] _RAND_2969;
  reg [31:0] _RAND_2970;
  reg [31:0] _RAND_2971;
  reg [31:0] _RAND_2972;
  reg [31:0] _RAND_2973;
  reg [31:0] _RAND_2974;
  reg [31:0] _RAND_2975;
  reg [31:0] _RAND_2976;
  reg [31:0] _RAND_2977;
  reg [31:0] _RAND_2978;
  reg [31:0] _RAND_2979;
  reg [31:0] _RAND_2980;
  reg [31:0] _RAND_2981;
  reg [31:0] _RAND_2982;
  reg [31:0] _RAND_2983;
  reg [31:0] _RAND_2984;
  reg [31:0] _RAND_2985;
  reg [31:0] _RAND_2986;
  reg [31:0] _RAND_2987;
  reg [31:0] _RAND_2988;
  reg [31:0] _RAND_2989;
  reg [31:0] _RAND_2990;
  reg [31:0] _RAND_2991;
  reg [31:0] _RAND_2992;
  reg [31:0] _RAND_2993;
  reg [31:0] _RAND_2994;
  reg [31:0] _RAND_2995;
  reg [31:0] _RAND_2996;
  reg [31:0] _RAND_2997;
  reg [31:0] _RAND_2998;
  reg [31:0] _RAND_2999;
  reg [31:0] _RAND_3000;
  reg [31:0] _RAND_3001;
  reg [31:0] _RAND_3002;
  reg [31:0] _RAND_3003;
  reg [31:0] _RAND_3004;
  reg [31:0] _RAND_3005;
  reg [31:0] _RAND_3006;
  reg [31:0] _RAND_3007;
  reg [31:0] _RAND_3008;
  reg [31:0] _RAND_3009;
  reg [31:0] _RAND_3010;
  reg [31:0] _RAND_3011;
  reg [31:0] _RAND_3012;
  reg [31:0] _RAND_3013;
  reg [31:0] _RAND_3014;
  reg [31:0] _RAND_3015;
  reg [31:0] _RAND_3016;
  reg [31:0] _RAND_3017;
  reg [31:0] _RAND_3018;
  reg [31:0] _RAND_3019;
  reg [31:0] _RAND_3020;
  reg [31:0] _RAND_3021;
  reg [31:0] _RAND_3022;
  reg [31:0] _RAND_3023;
  reg [31:0] _RAND_3024;
  reg [31:0] _RAND_3025;
  reg [31:0] _RAND_3026;
  reg [31:0] _RAND_3027;
  reg [31:0] _RAND_3028;
  reg [31:0] _RAND_3029;
  reg [31:0] _RAND_3030;
  reg [31:0] _RAND_3031;
  reg [31:0] _RAND_3032;
  reg [31:0] _RAND_3033;
  reg [31:0] _RAND_3034;
  reg [31:0] _RAND_3035;
  reg [31:0] _RAND_3036;
  reg [31:0] _RAND_3037;
  reg [31:0] _RAND_3038;
  reg [31:0] _RAND_3039;
  reg [31:0] _RAND_3040;
  reg [31:0] _RAND_3041;
  reg [31:0] _RAND_3042;
  reg [31:0] _RAND_3043;
  reg [31:0] _RAND_3044;
  reg [31:0] _RAND_3045;
  reg [31:0] _RAND_3046;
  reg [31:0] _RAND_3047;
  reg [31:0] _RAND_3048;
  reg [31:0] _RAND_3049;
  reg [31:0] _RAND_3050;
  reg [31:0] _RAND_3051;
  reg [31:0] _RAND_3052;
  reg [31:0] _RAND_3053;
  reg [31:0] _RAND_3054;
  reg [31:0] _RAND_3055;
  reg [31:0] _RAND_3056;
  reg [31:0] _RAND_3057;
  reg [31:0] _RAND_3058;
  reg [31:0] _RAND_3059;
  reg [31:0] _RAND_3060;
  reg [31:0] _RAND_3061;
  reg [31:0] _RAND_3062;
  reg [31:0] _RAND_3063;
  reg [31:0] _RAND_3064;
  reg [31:0] _RAND_3065;
  reg [31:0] _RAND_3066;
  reg [31:0] _RAND_3067;
  reg [31:0] _RAND_3068;
  reg [31:0] _RAND_3069;
  reg [31:0] _RAND_3070;
  reg [31:0] _RAND_3071;
  reg [31:0] _RAND_3072;
  reg [31:0] _RAND_3073;
  reg [31:0] _RAND_3074;
  reg [31:0] _RAND_3075;
  reg [31:0] _RAND_3076;
  reg [31:0] _RAND_3077;
  reg [31:0] _RAND_3078;
  reg [31:0] _RAND_3079;
  reg [31:0] _RAND_3080;
  reg [31:0] _RAND_3081;
  reg [31:0] _RAND_3082;
  reg [31:0] _RAND_3083;
  reg [31:0] _RAND_3084;
  reg [31:0] _RAND_3085;
  reg [31:0] _RAND_3086;
  reg [31:0] _RAND_3087;
  reg [31:0] _RAND_3088;
  reg [31:0] _RAND_3089;
  reg [31:0] _RAND_3090;
  reg [31:0] _RAND_3091;
  reg [31:0] _RAND_3092;
  reg [31:0] _RAND_3093;
  reg [31:0] _RAND_3094;
  reg [31:0] _RAND_3095;
  reg [31:0] _RAND_3096;
  reg [31:0] _RAND_3097;
  reg [31:0] _RAND_3098;
  reg [31:0] _RAND_3099;
  reg [31:0] _RAND_3100;
  reg [31:0] _RAND_3101;
  reg [31:0] _RAND_3102;
  reg [31:0] _RAND_3103;
  reg [31:0] _RAND_3104;
  reg [31:0] _RAND_3105;
  reg [31:0] _RAND_3106;
  reg [31:0] _RAND_3107;
  reg [31:0] _RAND_3108;
  reg [31:0] _RAND_3109;
  reg [31:0] _RAND_3110;
  reg [31:0] _RAND_3111;
  reg [31:0] _RAND_3112;
  reg [31:0] _RAND_3113;
  reg [31:0] _RAND_3114;
  reg [31:0] _RAND_3115;
  reg [31:0] _RAND_3116;
  reg [31:0] _RAND_3117;
  reg [31:0] _RAND_3118;
  reg [31:0] _RAND_3119;
  reg [31:0] _RAND_3120;
  reg [31:0] _RAND_3121;
  reg [31:0] _RAND_3122;
  reg [31:0] _RAND_3123;
  reg [31:0] _RAND_3124;
  reg [31:0] _RAND_3125;
  reg [31:0] _RAND_3126;
  reg [31:0] _RAND_3127;
  reg [31:0] _RAND_3128;
  reg [31:0] _RAND_3129;
  reg [31:0] _RAND_3130;
  reg [31:0] _RAND_3131;
  reg [31:0] _RAND_3132;
  reg [31:0] _RAND_3133;
  reg [31:0] _RAND_3134;
  reg [31:0] _RAND_3135;
  reg [31:0] _RAND_3136;
  reg [31:0] _RAND_3137;
  reg [31:0] _RAND_3138;
  reg [31:0] _RAND_3139;
  reg [31:0] _RAND_3140;
  reg [31:0] _RAND_3141;
  reg [31:0] _RAND_3142;
  reg [31:0] _RAND_3143;
  reg [31:0] _RAND_3144;
  reg [31:0] _RAND_3145;
  reg [31:0] _RAND_3146;
  reg [31:0] _RAND_3147;
  reg [31:0] _RAND_3148;
  reg [31:0] _RAND_3149;
  reg [31:0] _RAND_3150;
  reg [31:0] _RAND_3151;
  reg [31:0] _RAND_3152;
  reg [31:0] _RAND_3153;
  reg [31:0] _RAND_3154;
  reg [31:0] _RAND_3155;
  reg [31:0] _RAND_3156;
  reg [31:0] _RAND_3157;
  reg [31:0] _RAND_3158;
  reg [31:0] _RAND_3159;
  reg [31:0] _RAND_3160;
  reg [31:0] _RAND_3161;
  reg [31:0] _RAND_3162;
  reg [31:0] _RAND_3163;
  reg [31:0] _RAND_3164;
  reg [31:0] _RAND_3165;
  reg [31:0] _RAND_3166;
  reg [31:0] _RAND_3167;
  reg [31:0] _RAND_3168;
  reg [31:0] _RAND_3169;
  reg [31:0] _RAND_3170;
  reg [31:0] _RAND_3171;
  reg [31:0] _RAND_3172;
  reg [31:0] _RAND_3173;
  reg [31:0] _RAND_3174;
  reg [31:0] _RAND_3175;
  reg [31:0] _RAND_3176;
  reg [31:0] _RAND_3177;
  reg [31:0] _RAND_3178;
  reg [31:0] _RAND_3179;
  reg [31:0] _RAND_3180;
  reg [31:0] _RAND_3181;
  reg [31:0] _RAND_3182;
  reg [31:0] _RAND_3183;
  reg [31:0] _RAND_3184;
  reg [31:0] _RAND_3185;
  reg [31:0] _RAND_3186;
  reg [31:0] _RAND_3187;
  reg [31:0] _RAND_3188;
  reg [31:0] _RAND_3189;
  reg [31:0] _RAND_3190;
  reg [31:0] _RAND_3191;
  reg [31:0] _RAND_3192;
  reg [31:0] _RAND_3193;
  reg [31:0] _RAND_3194;
  reg [31:0] _RAND_3195;
  reg [31:0] _RAND_3196;
  reg [31:0] _RAND_3197;
  reg [31:0] _RAND_3198;
  reg [31:0] _RAND_3199;
  reg [31:0] _RAND_3200;
  reg [31:0] _RAND_3201;
  reg [31:0] _RAND_3202;
  reg [31:0] _RAND_3203;
  reg [31:0] _RAND_3204;
  reg [31:0] _RAND_3205;
  reg [31:0] _RAND_3206;
  reg [31:0] _RAND_3207;
  reg [31:0] _RAND_3208;
  reg [31:0] _RAND_3209;
  reg [31:0] _RAND_3210;
  reg [31:0] _RAND_3211;
  reg [31:0] _RAND_3212;
  reg [31:0] _RAND_3213;
  reg [31:0] _RAND_3214;
  reg [31:0] _RAND_3215;
  reg [31:0] _RAND_3216;
  reg [31:0] _RAND_3217;
  reg [31:0] _RAND_3218;
  reg [31:0] _RAND_3219;
  reg [31:0] _RAND_3220;
  reg [31:0] _RAND_3221;
  reg [31:0] _RAND_3222;
  reg [31:0] _RAND_3223;
  reg [31:0] _RAND_3224;
  reg [31:0] _RAND_3225;
  reg [31:0] _RAND_3226;
  reg [31:0] _RAND_3227;
  reg [31:0] _RAND_3228;
  reg [31:0] _RAND_3229;
  reg [31:0] _RAND_3230;
  reg [31:0] _RAND_3231;
  reg [31:0] _RAND_3232;
  reg [31:0] _RAND_3233;
  reg [31:0] _RAND_3234;
  reg [31:0] _RAND_3235;
  reg [31:0] _RAND_3236;
  reg [31:0] _RAND_3237;
  reg [31:0] _RAND_3238;
  reg [31:0] _RAND_3239;
  reg [31:0] _RAND_3240;
  reg [31:0] _RAND_3241;
  reg [31:0] _RAND_3242;
  reg [31:0] _RAND_3243;
  reg [31:0] _RAND_3244;
  reg [31:0] _RAND_3245;
  reg [31:0] _RAND_3246;
  reg [31:0] _RAND_3247;
  reg [31:0] _RAND_3248;
  reg [31:0] _RAND_3249;
  reg [31:0] _RAND_3250;
  reg [31:0] _RAND_3251;
  reg [31:0] _RAND_3252;
  reg [31:0] _RAND_3253;
  reg [31:0] _RAND_3254;
  reg [31:0] _RAND_3255;
  reg [31:0] _RAND_3256;
  reg [31:0] _RAND_3257;
  reg [31:0] _RAND_3258;
  reg [31:0] _RAND_3259;
  reg [31:0] _RAND_3260;
  reg [31:0] _RAND_3261;
  reg [31:0] _RAND_3262;
  reg [31:0] _RAND_3263;
  reg [31:0] _RAND_3264;
  reg [31:0] _RAND_3265;
  reg [31:0] _RAND_3266;
  reg [31:0] _RAND_3267;
  reg [31:0] _RAND_3268;
  reg [31:0] _RAND_3269;
  reg [31:0] _RAND_3270;
  reg [31:0] _RAND_3271;
  reg [31:0] _RAND_3272;
  reg [31:0] _RAND_3273;
  reg [31:0] _RAND_3274;
  reg [31:0] _RAND_3275;
  reg [31:0] _RAND_3276;
  reg [31:0] _RAND_3277;
  reg [31:0] _RAND_3278;
  reg [31:0] _RAND_3279;
  reg [31:0] _RAND_3280;
  reg [31:0] _RAND_3281;
  reg [31:0] _RAND_3282;
  reg [31:0] _RAND_3283;
  reg [31:0] _RAND_3284;
  reg [31:0] _RAND_3285;
  reg [31:0] _RAND_3286;
  reg [31:0] _RAND_3287;
  reg [31:0] _RAND_3288;
  reg [31:0] _RAND_3289;
  reg [31:0] _RAND_3290;
  reg [31:0] _RAND_3291;
  reg [31:0] _RAND_3292;
  reg [31:0] _RAND_3293;
  reg [31:0] _RAND_3294;
  reg [31:0] _RAND_3295;
  reg [31:0] _RAND_3296;
  reg [31:0] _RAND_3297;
  reg [31:0] _RAND_3298;
  reg [31:0] _RAND_3299;
  reg [31:0] _RAND_3300;
  reg [31:0] _RAND_3301;
  reg [31:0] _RAND_3302;
  reg [31:0] _RAND_3303;
  reg [31:0] _RAND_3304;
  reg [31:0] _RAND_3305;
  reg [31:0] _RAND_3306;
  reg [31:0] _RAND_3307;
  reg [31:0] _RAND_3308;
  reg [31:0] _RAND_3309;
  reg [31:0] _RAND_3310;
  reg [31:0] _RAND_3311;
  reg [31:0] _RAND_3312;
  reg [31:0] _RAND_3313;
  reg [31:0] _RAND_3314;
  reg [31:0] _RAND_3315;
  reg [31:0] _RAND_3316;
  reg [31:0] _RAND_3317;
  reg [31:0] _RAND_3318;
  reg [31:0] _RAND_3319;
  reg [31:0] _RAND_3320;
  reg [31:0] _RAND_3321;
  reg [31:0] _RAND_3322;
  reg [31:0] _RAND_3323;
  reg [31:0] _RAND_3324;
  reg [31:0] _RAND_3325;
  reg [31:0] _RAND_3326;
  reg [31:0] _RAND_3327;
  reg [31:0] _RAND_3328;
  reg [31:0] _RAND_3329;
  reg [31:0] _RAND_3330;
  reg [31:0] _RAND_3331;
  reg [31:0] _RAND_3332;
  reg [31:0] _RAND_3333;
  reg [31:0] _RAND_3334;
  reg [31:0] _RAND_3335;
  reg [31:0] _RAND_3336;
  reg [31:0] _RAND_3337;
  reg [31:0] _RAND_3338;
  reg [31:0] _RAND_3339;
  reg [31:0] _RAND_3340;
  reg [31:0] _RAND_3341;
  reg [31:0] _RAND_3342;
  reg [31:0] _RAND_3343;
  reg [31:0] _RAND_3344;
  reg [31:0] _RAND_3345;
  reg [31:0] _RAND_3346;
  reg [31:0] _RAND_3347;
  reg [31:0] _RAND_3348;
  reg [31:0] _RAND_3349;
  reg [31:0] _RAND_3350;
  reg [31:0] _RAND_3351;
  reg [31:0] _RAND_3352;
  reg [31:0] _RAND_3353;
  reg [31:0] _RAND_3354;
  reg [31:0] _RAND_3355;
  reg [31:0] _RAND_3356;
  reg [31:0] _RAND_3357;
  reg [31:0] _RAND_3358;
  reg [31:0] _RAND_3359;
  reg [31:0] _RAND_3360;
  reg [31:0] _RAND_3361;
  reg [31:0] _RAND_3362;
  reg [31:0] _RAND_3363;
  reg [31:0] _RAND_3364;
  reg [31:0] _RAND_3365;
  reg [31:0] _RAND_3366;
  reg [31:0] _RAND_3367;
  reg [31:0] _RAND_3368;
  reg [31:0] _RAND_3369;
  reg [31:0] _RAND_3370;
  reg [31:0] _RAND_3371;
  reg [31:0] _RAND_3372;
  reg [31:0] _RAND_3373;
  reg [31:0] _RAND_3374;
  reg [31:0] _RAND_3375;
  reg [31:0] _RAND_3376;
  reg [31:0] _RAND_3377;
  reg [31:0] _RAND_3378;
  reg [31:0] _RAND_3379;
  reg [31:0] _RAND_3380;
  reg [31:0] _RAND_3381;
  reg [31:0] _RAND_3382;
  reg [31:0] _RAND_3383;
  reg [31:0] _RAND_3384;
  reg [31:0] _RAND_3385;
  reg [31:0] _RAND_3386;
  reg [31:0] _RAND_3387;
  reg [31:0] _RAND_3388;
  reg [31:0] _RAND_3389;
  reg [31:0] _RAND_3390;
  reg [31:0] _RAND_3391;
  reg [31:0] _RAND_3392;
  reg [31:0] _RAND_3393;
  reg [31:0] _RAND_3394;
  reg [31:0] _RAND_3395;
  reg [31:0] _RAND_3396;
  reg [31:0] _RAND_3397;
  reg [31:0] _RAND_3398;
  reg [31:0] _RAND_3399;
  reg [31:0] _RAND_3400;
  reg [31:0] _RAND_3401;
  reg [31:0] _RAND_3402;
  reg [31:0] _RAND_3403;
  reg [31:0] _RAND_3404;
  reg [31:0] _RAND_3405;
  reg [31:0] _RAND_3406;
  reg [31:0] _RAND_3407;
  reg [31:0] _RAND_3408;
  reg [31:0] _RAND_3409;
  reg [31:0] _RAND_3410;
  reg [31:0] _RAND_3411;
  reg [31:0] _RAND_3412;
  reg [31:0] _RAND_3413;
  reg [31:0] _RAND_3414;
  reg [31:0] _RAND_3415;
  reg [31:0] _RAND_3416;
  reg [31:0] _RAND_3417;
  reg [31:0] _RAND_3418;
  reg [31:0] _RAND_3419;
  reg [31:0] _RAND_3420;
  reg [31:0] _RAND_3421;
  reg [31:0] _RAND_3422;
  reg [31:0] _RAND_3423;
  reg [31:0] _RAND_3424;
  reg [31:0] _RAND_3425;
  reg [31:0] _RAND_3426;
  reg [31:0] _RAND_3427;
  reg [31:0] _RAND_3428;
  reg [31:0] _RAND_3429;
  reg [31:0] _RAND_3430;
  reg [31:0] _RAND_3431;
  reg [31:0] _RAND_3432;
  reg [31:0] _RAND_3433;
  reg [31:0] _RAND_3434;
  reg [31:0] _RAND_3435;
  reg [31:0] _RAND_3436;
  reg [31:0] _RAND_3437;
  reg [31:0] _RAND_3438;
  reg [31:0] _RAND_3439;
  reg [31:0] _RAND_3440;
  reg [31:0] _RAND_3441;
  reg [31:0] _RAND_3442;
  reg [31:0] _RAND_3443;
  reg [31:0] _RAND_3444;
  reg [31:0] _RAND_3445;
  reg [31:0] _RAND_3446;
  reg [31:0] _RAND_3447;
  reg [31:0] _RAND_3448;
  reg [31:0] _RAND_3449;
  reg [31:0] _RAND_3450;
  reg [31:0] _RAND_3451;
  reg [31:0] _RAND_3452;
  reg [31:0] _RAND_3453;
  reg [31:0] _RAND_3454;
  reg [31:0] _RAND_3455;
  reg [31:0] _RAND_3456;
  reg [31:0] _RAND_3457;
  reg [31:0] _RAND_3458;
  reg [31:0] _RAND_3459;
  reg [31:0] _RAND_3460;
  reg [31:0] _RAND_3461;
  reg [31:0] _RAND_3462;
  reg [31:0] _RAND_3463;
  reg [31:0] _RAND_3464;
  reg [31:0] _RAND_3465;
  reg [31:0] _RAND_3466;
  reg [31:0] _RAND_3467;
  reg [31:0] _RAND_3468;
  reg [31:0] _RAND_3469;
  reg [31:0] _RAND_3470;
  reg [31:0] _RAND_3471;
  reg [31:0] _RAND_3472;
  reg [31:0] _RAND_3473;
  reg [31:0] _RAND_3474;
  reg [31:0] _RAND_3475;
  reg [31:0] _RAND_3476;
  reg [31:0] _RAND_3477;
  reg [31:0] _RAND_3478;
  reg [31:0] _RAND_3479;
  reg [31:0] _RAND_3480;
  reg [31:0] _RAND_3481;
  reg [31:0] _RAND_3482;
  reg [31:0] _RAND_3483;
  reg [31:0] _RAND_3484;
  reg [31:0] _RAND_3485;
  reg [31:0] _RAND_3486;
  reg [31:0] _RAND_3487;
  reg [31:0] _RAND_3488;
  reg [31:0] _RAND_3489;
  reg [31:0] _RAND_3490;
  reg [31:0] _RAND_3491;
  reg [31:0] _RAND_3492;
  reg [31:0] _RAND_3493;
  reg [31:0] _RAND_3494;
  reg [31:0] _RAND_3495;
  reg [31:0] _RAND_3496;
  reg [31:0] _RAND_3497;
  reg [31:0] _RAND_3498;
  reg [31:0] _RAND_3499;
  reg [31:0] _RAND_3500;
  reg [31:0] _RAND_3501;
  reg [31:0] _RAND_3502;
  reg [31:0] _RAND_3503;
  reg [31:0] _RAND_3504;
  reg [31:0] _RAND_3505;
  reg [31:0] _RAND_3506;
  reg [31:0] _RAND_3507;
  reg [31:0] _RAND_3508;
  reg [31:0] _RAND_3509;
  reg [31:0] _RAND_3510;
  reg [31:0] _RAND_3511;
  reg [31:0] _RAND_3512;
  reg [31:0] _RAND_3513;
  reg [31:0] _RAND_3514;
  reg [31:0] _RAND_3515;
  reg [31:0] _RAND_3516;
  reg [31:0] _RAND_3517;
  reg [31:0] _RAND_3518;
  reg [31:0] _RAND_3519;
  reg [31:0] _RAND_3520;
  reg [31:0] _RAND_3521;
  reg [31:0] _RAND_3522;
  reg [31:0] _RAND_3523;
  reg [31:0] _RAND_3524;
  reg [31:0] _RAND_3525;
  reg [31:0] _RAND_3526;
  reg [31:0] _RAND_3527;
  reg [31:0] _RAND_3528;
  reg [31:0] _RAND_3529;
  reg [31:0] _RAND_3530;
  reg [31:0] _RAND_3531;
  reg [31:0] _RAND_3532;
  reg [31:0] _RAND_3533;
  reg [31:0] _RAND_3534;
  reg [31:0] _RAND_3535;
  reg [31:0] _RAND_3536;
  reg [31:0] _RAND_3537;
  reg [31:0] _RAND_3538;
  reg [31:0] _RAND_3539;
  reg [31:0] _RAND_3540;
  reg [31:0] _RAND_3541;
  reg [31:0] _RAND_3542;
  reg [31:0] _RAND_3543;
  reg [31:0] _RAND_3544;
  reg [31:0] _RAND_3545;
  reg [31:0] _RAND_3546;
  reg [31:0] _RAND_3547;
  reg [31:0] _RAND_3548;
  reg [31:0] _RAND_3549;
  reg [31:0] _RAND_3550;
  reg [31:0] _RAND_3551;
  reg [31:0] _RAND_3552;
  reg [31:0] _RAND_3553;
  reg [31:0] _RAND_3554;
  reg [31:0] _RAND_3555;
  reg [31:0] _RAND_3556;
  reg [31:0] _RAND_3557;
  reg [31:0] _RAND_3558;
  reg [31:0] _RAND_3559;
  reg [31:0] _RAND_3560;
  reg [31:0] _RAND_3561;
  reg [31:0] _RAND_3562;
  reg [31:0] _RAND_3563;
  reg [31:0] _RAND_3564;
  reg [31:0] _RAND_3565;
  reg [31:0] _RAND_3566;
  reg [31:0] _RAND_3567;
  reg [31:0] _RAND_3568;
  reg [31:0] _RAND_3569;
  reg [31:0] _RAND_3570;
  reg [31:0] _RAND_3571;
  reg [31:0] _RAND_3572;
  reg [31:0] _RAND_3573;
  reg [31:0] _RAND_3574;
  reg [31:0] _RAND_3575;
  reg [31:0] _RAND_3576;
  reg [31:0] _RAND_3577;
  reg [31:0] _RAND_3578;
  reg [31:0] _RAND_3579;
  reg [31:0] _RAND_3580;
  reg [31:0] _RAND_3581;
  reg [31:0] _RAND_3582;
  reg [31:0] _RAND_3583;
  reg [31:0] _RAND_3584;
  reg [31:0] _RAND_3585;
  reg [31:0] _RAND_3586;
  reg [31:0] _RAND_3587;
  reg [31:0] _RAND_3588;
  reg [31:0] _RAND_3589;
  reg [31:0] _RAND_3590;
  reg [31:0] _RAND_3591;
  reg [31:0] _RAND_3592;
  reg [31:0] _RAND_3593;
  reg [31:0] _RAND_3594;
  reg [31:0] _RAND_3595;
  reg [31:0] _RAND_3596;
  reg [31:0] _RAND_3597;
  reg [31:0] _RAND_3598;
  reg [31:0] _RAND_3599;
  reg [31:0] _RAND_3600;
  reg [31:0] _RAND_3601;
  reg [31:0] _RAND_3602;
  reg [31:0] _RAND_3603;
  reg [31:0] _RAND_3604;
  reg [31:0] _RAND_3605;
  reg [31:0] _RAND_3606;
  reg [31:0] _RAND_3607;
  reg [31:0] _RAND_3608;
  reg [31:0] _RAND_3609;
  reg [31:0] _RAND_3610;
  reg [31:0] _RAND_3611;
  reg [31:0] _RAND_3612;
  reg [31:0] _RAND_3613;
  reg [31:0] _RAND_3614;
  reg [31:0] _RAND_3615;
  reg [31:0] _RAND_3616;
  reg [31:0] _RAND_3617;
  reg [31:0] _RAND_3618;
  reg [31:0] _RAND_3619;
  reg [31:0] _RAND_3620;
  reg [31:0] _RAND_3621;
  reg [31:0] _RAND_3622;
  reg [31:0] _RAND_3623;
  reg [31:0] _RAND_3624;
  reg [31:0] _RAND_3625;
  reg [31:0] _RAND_3626;
  reg [31:0] _RAND_3627;
  reg [31:0] _RAND_3628;
  reg [31:0] _RAND_3629;
  reg [31:0] _RAND_3630;
  reg [31:0] _RAND_3631;
  reg [31:0] _RAND_3632;
  reg [31:0] _RAND_3633;
  reg [31:0] _RAND_3634;
  reg [31:0] _RAND_3635;
  reg [31:0] _RAND_3636;
  reg [31:0] _RAND_3637;
  reg [31:0] _RAND_3638;
  reg [31:0] _RAND_3639;
  reg [31:0] _RAND_3640;
  reg [31:0] _RAND_3641;
  reg [31:0] _RAND_3642;
  reg [31:0] _RAND_3643;
  reg [31:0] _RAND_3644;
  reg [31:0] _RAND_3645;
  reg [31:0] _RAND_3646;
  reg [31:0] _RAND_3647;
  reg [31:0] _RAND_3648;
  reg [31:0] _RAND_3649;
  reg [31:0] _RAND_3650;
  reg [31:0] _RAND_3651;
  reg [31:0] _RAND_3652;
  reg [31:0] _RAND_3653;
  reg [31:0] _RAND_3654;
  reg [31:0] _RAND_3655;
  reg [31:0] _RAND_3656;
  reg [31:0] _RAND_3657;
  reg [31:0] _RAND_3658;
  reg [31:0] _RAND_3659;
  reg [31:0] _RAND_3660;
  reg [31:0] _RAND_3661;
  reg [31:0] _RAND_3662;
  reg [31:0] _RAND_3663;
  reg [31:0] _RAND_3664;
  reg [31:0] _RAND_3665;
  reg [31:0] _RAND_3666;
  reg [31:0] _RAND_3667;
  reg [31:0] _RAND_3668;
  reg [31:0] _RAND_3669;
  reg [31:0] _RAND_3670;
  reg [31:0] _RAND_3671;
  reg [31:0] _RAND_3672;
  reg [31:0] _RAND_3673;
  reg [31:0] _RAND_3674;
  reg [31:0] _RAND_3675;
  reg [31:0] _RAND_3676;
  reg [31:0] _RAND_3677;
  reg [31:0] _RAND_3678;
  reg [31:0] _RAND_3679;
  reg [31:0] _RAND_3680;
  reg [31:0] _RAND_3681;
  reg [31:0] _RAND_3682;
  reg [31:0] _RAND_3683;
  reg [31:0] _RAND_3684;
  reg [31:0] _RAND_3685;
  reg [31:0] _RAND_3686;
  reg [31:0] _RAND_3687;
  reg [31:0] _RAND_3688;
  reg [31:0] _RAND_3689;
  reg [31:0] _RAND_3690;
  reg [31:0] _RAND_3691;
  reg [31:0] _RAND_3692;
  reg [31:0] _RAND_3693;
  reg [31:0] _RAND_3694;
  reg [31:0] _RAND_3695;
  reg [31:0] _RAND_3696;
  reg [31:0] _RAND_3697;
  reg [31:0] _RAND_3698;
  reg [31:0] _RAND_3699;
  reg [31:0] _RAND_3700;
  reg [31:0] _RAND_3701;
  reg [31:0] _RAND_3702;
  reg [31:0] _RAND_3703;
  reg [31:0] _RAND_3704;
  reg [31:0] _RAND_3705;
  reg [31:0] _RAND_3706;
  reg [31:0] _RAND_3707;
  reg [31:0] _RAND_3708;
  reg [31:0] _RAND_3709;
  reg [31:0] _RAND_3710;
  reg [31:0] _RAND_3711;
  reg [31:0] _RAND_3712;
  reg [31:0] _RAND_3713;
  reg [31:0] _RAND_3714;
  reg [31:0] _RAND_3715;
  reg [31:0] _RAND_3716;
  reg [31:0] _RAND_3717;
  reg [31:0] _RAND_3718;
  reg [31:0] _RAND_3719;
  reg [31:0] _RAND_3720;
  reg [31:0] _RAND_3721;
  reg [31:0] _RAND_3722;
  reg [31:0] _RAND_3723;
  reg [31:0] _RAND_3724;
  reg [31:0] _RAND_3725;
  reg [31:0] _RAND_3726;
  reg [31:0] _RAND_3727;
  reg [31:0] _RAND_3728;
  reg [31:0] _RAND_3729;
  reg [31:0] _RAND_3730;
  reg [31:0] _RAND_3731;
  reg [31:0] _RAND_3732;
  reg [31:0] _RAND_3733;
  reg [31:0] _RAND_3734;
  reg [31:0] _RAND_3735;
  reg [31:0] _RAND_3736;
  reg [31:0] _RAND_3737;
  reg [31:0] _RAND_3738;
  reg [31:0] _RAND_3739;
  reg [31:0] _RAND_3740;
  reg [31:0] _RAND_3741;
  reg [31:0] _RAND_3742;
  reg [31:0] _RAND_3743;
  reg [31:0] _RAND_3744;
  reg [31:0] _RAND_3745;
  reg [31:0] _RAND_3746;
  reg [31:0] _RAND_3747;
  reg [31:0] _RAND_3748;
  reg [31:0] _RAND_3749;
  reg [31:0] _RAND_3750;
  reg [31:0] _RAND_3751;
  reg [31:0] _RAND_3752;
  reg [31:0] _RAND_3753;
  reg [31:0] _RAND_3754;
  reg [31:0] _RAND_3755;
  reg [31:0] _RAND_3756;
  reg [31:0] _RAND_3757;
  reg [31:0] _RAND_3758;
  reg [31:0] _RAND_3759;
  reg [31:0] _RAND_3760;
  reg [31:0] _RAND_3761;
  reg [31:0] _RAND_3762;
  reg [31:0] _RAND_3763;
  reg [31:0] _RAND_3764;
  reg [31:0] _RAND_3765;
  reg [31:0] _RAND_3766;
  reg [31:0] _RAND_3767;
  reg [31:0] _RAND_3768;
  reg [31:0] _RAND_3769;
  reg [31:0] _RAND_3770;
  reg [31:0] _RAND_3771;
  reg [31:0] _RAND_3772;
  reg [31:0] _RAND_3773;
  reg [31:0] _RAND_3774;
  reg [31:0] _RAND_3775;
  reg [31:0] _RAND_3776;
  reg [31:0] _RAND_3777;
  reg [31:0] _RAND_3778;
  reg [31:0] _RAND_3779;
  reg [31:0] _RAND_3780;
  reg [31:0] _RAND_3781;
  reg [31:0] _RAND_3782;
  reg [31:0] _RAND_3783;
  reg [31:0] _RAND_3784;
  reg [31:0] _RAND_3785;
  reg [31:0] _RAND_3786;
  reg [31:0] _RAND_3787;
  reg [31:0] _RAND_3788;
  reg [31:0] _RAND_3789;
  reg [31:0] _RAND_3790;
  reg [31:0] _RAND_3791;
  reg [31:0] _RAND_3792;
  reg [31:0] _RAND_3793;
  reg [31:0] _RAND_3794;
  reg [31:0] _RAND_3795;
  reg [31:0] _RAND_3796;
  reg [31:0] _RAND_3797;
  reg [31:0] _RAND_3798;
  reg [31:0] _RAND_3799;
  reg [31:0] _RAND_3800;
  reg [31:0] _RAND_3801;
  reg [31:0] _RAND_3802;
  reg [31:0] _RAND_3803;
  reg [31:0] _RAND_3804;
  reg [31:0] _RAND_3805;
  reg [31:0] _RAND_3806;
  reg [31:0] _RAND_3807;
  reg [31:0] _RAND_3808;
  reg [31:0] _RAND_3809;
  reg [31:0] _RAND_3810;
  reg [31:0] _RAND_3811;
  reg [31:0] _RAND_3812;
  reg [31:0] _RAND_3813;
  reg [31:0] _RAND_3814;
  reg [31:0] _RAND_3815;
  reg [31:0] _RAND_3816;
  reg [31:0] _RAND_3817;
  reg [31:0] _RAND_3818;
  reg [31:0] _RAND_3819;
  reg [31:0] _RAND_3820;
  reg [31:0] _RAND_3821;
  reg [31:0] _RAND_3822;
  reg [31:0] _RAND_3823;
  reg [31:0] _RAND_3824;
  reg [31:0] _RAND_3825;
  reg [31:0] _RAND_3826;
  reg [31:0] _RAND_3827;
  reg [31:0] _RAND_3828;
  reg [31:0] _RAND_3829;
  reg [31:0] _RAND_3830;
  reg [31:0] _RAND_3831;
  reg [31:0] _RAND_3832;
  reg [31:0] _RAND_3833;
  reg [31:0] _RAND_3834;
  reg [31:0] _RAND_3835;
  reg [31:0] _RAND_3836;
  reg [31:0] _RAND_3837;
  reg [31:0] _RAND_3838;
  reg [31:0] _RAND_3839;
  reg [31:0] _RAND_3840;
  reg [31:0] _RAND_3841;
  reg [31:0] _RAND_3842;
  reg [31:0] _RAND_3843;
  reg [31:0] _RAND_3844;
  reg [31:0] _RAND_3845;
  reg [31:0] _RAND_3846;
  reg [31:0] _RAND_3847;
  reg [31:0] _RAND_3848;
  reg [31:0] _RAND_3849;
  reg [31:0] _RAND_3850;
  reg [31:0] _RAND_3851;
  reg [31:0] _RAND_3852;
  reg [31:0] _RAND_3853;
  reg [31:0] _RAND_3854;
  reg [31:0] _RAND_3855;
  reg [31:0] _RAND_3856;
  reg [31:0] _RAND_3857;
  reg [31:0] _RAND_3858;
  reg [31:0] _RAND_3859;
  reg [31:0] _RAND_3860;
  reg [31:0] _RAND_3861;
  reg [31:0] _RAND_3862;
  reg [31:0] _RAND_3863;
  reg [31:0] _RAND_3864;
  reg [31:0] _RAND_3865;
  reg [31:0] _RAND_3866;
  reg [31:0] _RAND_3867;
  reg [31:0] _RAND_3868;
  reg [31:0] _RAND_3869;
  reg [31:0] _RAND_3870;
  reg [31:0] _RAND_3871;
  reg [31:0] _RAND_3872;
  reg [31:0] _RAND_3873;
  reg [31:0] _RAND_3874;
  reg [31:0] _RAND_3875;
  reg [31:0] _RAND_3876;
  reg [31:0] _RAND_3877;
  reg [31:0] _RAND_3878;
  reg [31:0] _RAND_3879;
  reg [31:0] _RAND_3880;
  reg [31:0] _RAND_3881;
  reg [31:0] _RAND_3882;
  reg [31:0] _RAND_3883;
  reg [31:0] _RAND_3884;
  reg [31:0] _RAND_3885;
  reg [31:0] _RAND_3886;
  reg [31:0] _RAND_3887;
  reg [31:0] _RAND_3888;
  reg [31:0] _RAND_3889;
  reg [31:0] _RAND_3890;
  reg [31:0] _RAND_3891;
  reg [31:0] _RAND_3892;
  reg [31:0] _RAND_3893;
  reg [31:0] _RAND_3894;
  reg [31:0] _RAND_3895;
  reg [31:0] _RAND_3896;
  reg [31:0] _RAND_3897;
  reg [31:0] _RAND_3898;
  reg [31:0] _RAND_3899;
  reg [31:0] _RAND_3900;
  reg [31:0] _RAND_3901;
  reg [31:0] _RAND_3902;
  reg [31:0] _RAND_3903;
  reg [31:0] _RAND_3904;
  reg [31:0] _RAND_3905;
  reg [31:0] _RAND_3906;
  reg [31:0] _RAND_3907;
  reg [31:0] _RAND_3908;
  reg [31:0] _RAND_3909;
  reg [31:0] _RAND_3910;
  reg [31:0] _RAND_3911;
  reg [31:0] _RAND_3912;
  reg [31:0] _RAND_3913;
  reg [31:0] _RAND_3914;
  reg [31:0] _RAND_3915;
  reg [31:0] _RAND_3916;
  reg [31:0] _RAND_3917;
  reg [31:0] _RAND_3918;
  reg [31:0] _RAND_3919;
  reg [31:0] _RAND_3920;
  reg [31:0] _RAND_3921;
  reg [31:0] _RAND_3922;
  reg [31:0] _RAND_3923;
  reg [31:0] _RAND_3924;
  reg [31:0] _RAND_3925;
  reg [31:0] _RAND_3926;
  reg [31:0] _RAND_3927;
  reg [31:0] _RAND_3928;
  reg [31:0] _RAND_3929;
  reg [31:0] _RAND_3930;
  reg [31:0] _RAND_3931;
  reg [31:0] _RAND_3932;
  reg [31:0] _RAND_3933;
  reg [31:0] _RAND_3934;
  reg [31:0] _RAND_3935;
  reg [31:0] _RAND_3936;
  reg [31:0] _RAND_3937;
  reg [31:0] _RAND_3938;
  reg [31:0] _RAND_3939;
  reg [31:0] _RAND_3940;
  reg [31:0] _RAND_3941;
  reg [31:0] _RAND_3942;
  reg [31:0] _RAND_3943;
  reg [31:0] _RAND_3944;
  reg [31:0] _RAND_3945;
  reg [31:0] _RAND_3946;
  reg [31:0] _RAND_3947;
  reg [31:0] _RAND_3948;
  reg [31:0] _RAND_3949;
  reg [31:0] _RAND_3950;
  reg [31:0] _RAND_3951;
  reg [31:0] _RAND_3952;
  reg [31:0] _RAND_3953;
  reg [31:0] _RAND_3954;
  reg [31:0] _RAND_3955;
  reg [31:0] _RAND_3956;
  reg [31:0] _RAND_3957;
  reg [31:0] _RAND_3958;
  reg [31:0] _RAND_3959;
  reg [31:0] _RAND_3960;
  reg [31:0] _RAND_3961;
  reg [31:0] _RAND_3962;
  reg [31:0] _RAND_3963;
  reg [31:0] _RAND_3964;
  reg [31:0] _RAND_3965;
  reg [31:0] _RAND_3966;
  reg [31:0] _RAND_3967;
  reg [31:0] _RAND_3968;
  reg [31:0] _RAND_3969;
  reg [31:0] _RAND_3970;
  reg [31:0] _RAND_3971;
  reg [31:0] _RAND_3972;
  reg [31:0] _RAND_3973;
  reg [31:0] _RAND_3974;
  reg [31:0] _RAND_3975;
  reg [31:0] _RAND_3976;
  reg [31:0] _RAND_3977;
  reg [31:0] _RAND_3978;
  reg [31:0] _RAND_3979;
  reg [31:0] _RAND_3980;
  reg [31:0] _RAND_3981;
  reg [31:0] _RAND_3982;
  reg [31:0] _RAND_3983;
  reg [31:0] _RAND_3984;
  reg [31:0] _RAND_3985;
  reg [31:0] _RAND_3986;
  reg [31:0] _RAND_3987;
  reg [31:0] _RAND_3988;
  reg [31:0] _RAND_3989;
  reg [31:0] _RAND_3990;
  reg [31:0] _RAND_3991;
  reg [31:0] _RAND_3992;
  reg [31:0] _RAND_3993;
  reg [31:0] _RAND_3994;
  reg [31:0] _RAND_3995;
  reg [31:0] _RAND_3996;
  reg [31:0] _RAND_3997;
  reg [31:0] _RAND_3998;
  reg [31:0] _RAND_3999;
  reg [31:0] _RAND_4000;
  reg [31:0] _RAND_4001;
  reg [31:0] _RAND_4002;
  reg [31:0] _RAND_4003;
  reg [31:0] _RAND_4004;
  reg [31:0] _RAND_4005;
  reg [31:0] _RAND_4006;
  reg [31:0] _RAND_4007;
  reg [31:0] _RAND_4008;
  reg [31:0] _RAND_4009;
  reg [31:0] _RAND_4010;
  reg [31:0] _RAND_4011;
  reg [31:0] _RAND_4012;
  reg [31:0] _RAND_4013;
  reg [31:0] _RAND_4014;
  reg [31:0] _RAND_4015;
  reg [31:0] _RAND_4016;
  reg [31:0] _RAND_4017;
  reg [31:0] _RAND_4018;
  reg [31:0] _RAND_4019;
  reg [31:0] _RAND_4020;
  reg [31:0] _RAND_4021;
  reg [31:0] _RAND_4022;
  reg [31:0] _RAND_4023;
  reg [31:0] _RAND_4024;
  reg [31:0] _RAND_4025;
  reg [31:0] _RAND_4026;
  reg [31:0] _RAND_4027;
  reg [31:0] _RAND_4028;
  reg [31:0] _RAND_4029;
  reg [31:0] _RAND_4030;
  reg [31:0] _RAND_4031;
  reg [31:0] _RAND_4032;
  reg [31:0] _RAND_4033;
  reg [31:0] _RAND_4034;
  reg [31:0] _RAND_4035;
  reg [31:0] _RAND_4036;
  reg [31:0] _RAND_4037;
  reg [31:0] _RAND_4038;
  reg [31:0] _RAND_4039;
  reg [31:0] _RAND_4040;
  reg [31:0] _RAND_4041;
  reg [31:0] _RAND_4042;
  reg [31:0] _RAND_4043;
  reg [31:0] _RAND_4044;
  reg [31:0] _RAND_4045;
  reg [31:0] _RAND_4046;
  reg [31:0] _RAND_4047;
  reg [31:0] _RAND_4048;
  reg [31:0] _RAND_4049;
  reg [31:0] _RAND_4050;
  reg [31:0] _RAND_4051;
  reg [31:0] _RAND_4052;
  reg [31:0] _RAND_4053;
  reg [31:0] _RAND_4054;
  reg [31:0] _RAND_4055;
  reg [31:0] _RAND_4056;
  reg [31:0] _RAND_4057;
  reg [31:0] _RAND_4058;
  reg [31:0] _RAND_4059;
  reg [31:0] _RAND_4060;
  reg [31:0] _RAND_4061;
  reg [31:0] _RAND_4062;
  reg [31:0] _RAND_4063;
  reg [31:0] _RAND_4064;
  reg [31:0] _RAND_4065;
  reg [31:0] _RAND_4066;
  reg [31:0] _RAND_4067;
  reg [31:0] _RAND_4068;
  reg [31:0] _RAND_4069;
  reg [31:0] _RAND_4070;
  reg [31:0] _RAND_4071;
  reg [31:0] _RAND_4072;
  reg [31:0] _RAND_4073;
  reg [31:0] _RAND_4074;
  reg [31:0] _RAND_4075;
  reg [31:0] _RAND_4076;
  reg [31:0] _RAND_4077;
  reg [31:0] _RAND_4078;
  reg [31:0] _RAND_4079;
  reg [31:0] _RAND_4080;
  reg [31:0] _RAND_4081;
  reg [31:0] _RAND_4082;
  reg [31:0] _RAND_4083;
  reg [31:0] _RAND_4084;
  reg [31:0] _RAND_4085;
  reg [31:0] _RAND_4086;
  reg [31:0] _RAND_4087;
  reg [31:0] _RAND_4088;
  reg [31:0] _RAND_4089;
  reg [31:0] _RAND_4090;
  reg [31:0] _RAND_4091;
  reg [31:0] _RAND_4092;
  reg [31:0] _RAND_4093;
  reg [31:0] _RAND_4094;
  reg [31:0] _RAND_4095;
  reg [31:0] _RAND_4096;
  reg [31:0] _RAND_4097;
  reg [31:0] _RAND_4098;
  reg [31:0] _RAND_4099;
  reg [31:0] _RAND_4100;
  reg [31:0] _RAND_4101;
  reg [31:0] _RAND_4102;
  reg [31:0] _RAND_4103;
  reg [31:0] _RAND_4104;
  reg [31:0] _RAND_4105;
  reg [31:0] _RAND_4106;
  reg [31:0] _RAND_4107;
  reg [31:0] _RAND_4108;
  reg [31:0] _RAND_4109;
  reg [31:0] _RAND_4110;
  reg [31:0] _RAND_4111;
  reg [31:0] _RAND_4112;
  reg [31:0] _RAND_4113;
  reg [31:0] _RAND_4114;
  reg [31:0] _RAND_4115;
  reg [31:0] _RAND_4116;
  reg [31:0] _RAND_4117;
  reg [31:0] _RAND_4118;
  reg [31:0] _RAND_4119;
  reg [31:0] _RAND_4120;
  reg [31:0] _RAND_4121;
  reg [31:0] _RAND_4122;
  reg [31:0] _RAND_4123;
  reg [31:0] _RAND_4124;
  reg [31:0] _RAND_4125;
  reg [31:0] _RAND_4126;
  reg [31:0] _RAND_4127;
  reg [31:0] _RAND_4128;
  reg [31:0] _RAND_4129;
  reg [31:0] _RAND_4130;
  reg [31:0] _RAND_4131;
  reg [31:0] _RAND_4132;
  reg [31:0] _RAND_4133;
  reg [31:0] _RAND_4134;
  reg [31:0] _RAND_4135;
  reg [31:0] _RAND_4136;
  reg [31:0] _RAND_4137;
  reg [31:0] _RAND_4138;
  reg [31:0] _RAND_4139;
  reg [31:0] _RAND_4140;
  reg [31:0] _RAND_4141;
  reg [31:0] _RAND_4142;
  reg [31:0] _RAND_4143;
  reg [31:0] _RAND_4144;
  reg [31:0] _RAND_4145;
  reg [31:0] _RAND_4146;
  reg [31:0] _RAND_4147;
  reg [31:0] _RAND_4148;
  reg [31:0] _RAND_4149;
  reg [31:0] _RAND_4150;
  reg [31:0] _RAND_4151;
  reg [31:0] _RAND_4152;
  reg [31:0] _RAND_4153;
  reg [31:0] _RAND_4154;
  reg [31:0] _RAND_4155;
  reg [31:0] _RAND_4156;
  reg [31:0] _RAND_4157;
  reg [31:0] _RAND_4158;
  reg [31:0] _RAND_4159;
  reg [31:0] _RAND_4160;
  reg [31:0] _RAND_4161;
  reg [31:0] _RAND_4162;
  reg [31:0] _RAND_4163;
  reg [31:0] _RAND_4164;
  reg [31:0] _RAND_4165;
  reg [31:0] _RAND_4166;
  reg [31:0] _RAND_4167;
  reg [31:0] _RAND_4168;
  reg [31:0] _RAND_4169;
  reg [31:0] _RAND_4170;
  reg [31:0] _RAND_4171;
  reg [31:0] _RAND_4172;
  reg [31:0] _RAND_4173;
  reg [31:0] _RAND_4174;
  reg [31:0] _RAND_4175;
  reg [31:0] _RAND_4176;
  reg [31:0] _RAND_4177;
  reg [31:0] _RAND_4178;
  reg [31:0] _RAND_4179;
  reg [31:0] _RAND_4180;
  reg [31:0] _RAND_4181;
  reg [31:0] _RAND_4182;
  reg [31:0] _RAND_4183;
  reg [31:0] _RAND_4184;
  reg [31:0] _RAND_4185;
  reg [31:0] _RAND_4186;
  reg [31:0] _RAND_4187;
  reg [31:0] _RAND_4188;
  reg [31:0] _RAND_4189;
  reg [31:0] _RAND_4190;
  reg [31:0] _RAND_4191;
  reg [31:0] _RAND_4192;
  reg [31:0] _RAND_4193;
  reg [31:0] _RAND_4194;
  reg [31:0] _RAND_4195;
  reg [31:0] _RAND_4196;
  reg [31:0] _RAND_4197;
  reg [31:0] _RAND_4198;
  reg [31:0] _RAND_4199;
  reg [31:0] _RAND_4200;
  reg [31:0] _RAND_4201;
  reg [31:0] _RAND_4202;
  reg [31:0] _RAND_4203;
  reg [31:0] _RAND_4204;
  reg [31:0] _RAND_4205;
  reg [31:0] _RAND_4206;
  reg [31:0] _RAND_4207;
  reg [31:0] _RAND_4208;
  reg [31:0] _RAND_4209;
  reg [31:0] _RAND_4210;
  reg [31:0] _RAND_4211;
  reg [31:0] _RAND_4212;
  reg [31:0] _RAND_4213;
  reg [31:0] _RAND_4214;
  reg [31:0] _RAND_4215;
  reg [31:0] _RAND_4216;
  reg [31:0] _RAND_4217;
  reg [31:0] _RAND_4218;
  reg [31:0] _RAND_4219;
  reg [31:0] _RAND_4220;
  reg [31:0] _RAND_4221;
  reg [31:0] _RAND_4222;
  reg [31:0] _RAND_4223;
  reg [31:0] _RAND_4224;
  reg [31:0] _RAND_4225;
  reg [31:0] _RAND_4226;
  reg [31:0] _RAND_4227;
  reg [31:0] _RAND_4228;
  reg [31:0] _RAND_4229;
  reg [31:0] _RAND_4230;
  reg [31:0] _RAND_4231;
  reg [31:0] _RAND_4232;
  reg [31:0] _RAND_4233;
  reg [31:0] _RAND_4234;
  reg [31:0] _RAND_4235;
  reg [31:0] _RAND_4236;
  reg [31:0] _RAND_4237;
  reg [31:0] _RAND_4238;
  reg [31:0] _RAND_4239;
  reg [31:0] _RAND_4240;
  reg [31:0] _RAND_4241;
  reg [31:0] _RAND_4242;
  reg [31:0] _RAND_4243;
  reg [31:0] _RAND_4244;
  reg [31:0] _RAND_4245;
  reg [31:0] _RAND_4246;
  reg [31:0] _RAND_4247;
  reg [31:0] _RAND_4248;
  reg [31:0] _RAND_4249;
  reg [31:0] _RAND_4250;
  reg [31:0] _RAND_4251;
  reg [31:0] _RAND_4252;
  reg [31:0] _RAND_4253;
  reg [31:0] _RAND_4254;
  reg [31:0] _RAND_4255;
  reg [31:0] _RAND_4256;
  reg [31:0] _RAND_4257;
  reg [31:0] _RAND_4258;
  reg [31:0] _RAND_4259;
  reg [31:0] _RAND_4260;
  reg [31:0] _RAND_4261;
  reg [31:0] _RAND_4262;
  reg [31:0] _RAND_4263;
  reg [31:0] _RAND_4264;
  reg [31:0] _RAND_4265;
  reg [31:0] _RAND_4266;
  reg [31:0] _RAND_4267;
  reg [31:0] _RAND_4268;
  reg [31:0] _RAND_4269;
  reg [31:0] _RAND_4270;
  reg [31:0] _RAND_4271;
  reg [31:0] _RAND_4272;
  reg [31:0] _RAND_4273;
  reg [31:0] _RAND_4274;
  reg [31:0] _RAND_4275;
  reg [31:0] _RAND_4276;
  reg [31:0] _RAND_4277;
  reg [31:0] _RAND_4278;
  reg [31:0] _RAND_4279;
  reg [31:0] _RAND_4280;
  reg [31:0] _RAND_4281;
  reg [31:0] _RAND_4282;
  reg [31:0] _RAND_4283;
  reg [31:0] _RAND_4284;
  reg [31:0] _RAND_4285;
  reg [31:0] _RAND_4286;
  reg [31:0] _RAND_4287;
  reg [31:0] _RAND_4288;
  reg [31:0] _RAND_4289;
  reg [31:0] _RAND_4290;
  reg [31:0] _RAND_4291;
  reg [31:0] _RAND_4292;
  reg [31:0] _RAND_4293;
  reg [31:0] _RAND_4294;
  reg [31:0] _RAND_4295;
  reg [31:0] _RAND_4296;
  reg [31:0] _RAND_4297;
  reg [31:0] _RAND_4298;
  reg [31:0] _RAND_4299;
  reg [31:0] _RAND_4300;
  reg [31:0] _RAND_4301;
  reg [31:0] _RAND_4302;
  reg [31:0] _RAND_4303;
  reg [31:0] _RAND_4304;
  reg [31:0] _RAND_4305;
  reg [31:0] _RAND_4306;
  reg [31:0] _RAND_4307;
  reg [31:0] _RAND_4308;
  reg [31:0] _RAND_4309;
  reg [31:0] _RAND_4310;
  reg [31:0] _RAND_4311;
  reg [31:0] _RAND_4312;
  reg [31:0] _RAND_4313;
  reg [31:0] _RAND_4314;
  reg [31:0] _RAND_4315;
  reg [31:0] _RAND_4316;
  reg [31:0] _RAND_4317;
  reg [31:0] _RAND_4318;
  reg [31:0] _RAND_4319;
  reg [31:0] _RAND_4320;
  reg [31:0] _RAND_4321;
  reg [31:0] _RAND_4322;
  reg [31:0] _RAND_4323;
  reg [31:0] _RAND_4324;
  reg [31:0] _RAND_4325;
  reg [31:0] _RAND_4326;
  reg [31:0] _RAND_4327;
  reg [31:0] _RAND_4328;
  reg [31:0] _RAND_4329;
  reg [31:0] _RAND_4330;
  reg [31:0] _RAND_4331;
  reg [31:0] _RAND_4332;
  reg [31:0] _RAND_4333;
  reg [31:0] _RAND_4334;
  reg [31:0] _RAND_4335;
  reg [31:0] _RAND_4336;
  reg [31:0] _RAND_4337;
  reg [31:0] _RAND_4338;
  reg [31:0] _RAND_4339;
  reg [31:0] _RAND_4340;
  reg [31:0] _RAND_4341;
  reg [31:0] _RAND_4342;
  reg [31:0] _RAND_4343;
  reg [31:0] _RAND_4344;
  reg [31:0] _RAND_4345;
  reg [31:0] _RAND_4346;
  reg [31:0] _RAND_4347;
  reg [31:0] _RAND_4348;
  reg [31:0] _RAND_4349;
  reg [31:0] _RAND_4350;
  reg [31:0] _RAND_4351;
  reg [31:0] _RAND_4352;
  reg [31:0] _RAND_4353;
  reg [31:0] _RAND_4354;
  reg [31:0] _RAND_4355;
  reg [31:0] _RAND_4356;
  reg [31:0] _RAND_4357;
  reg [31:0] _RAND_4358;
  reg [31:0] _RAND_4359;
  reg [31:0] _RAND_4360;
  reg [31:0] _RAND_4361;
  reg [31:0] _RAND_4362;
  reg [31:0] _RAND_4363;
  reg [31:0] _RAND_4364;
  reg [31:0] _RAND_4365;
  reg [31:0] _RAND_4366;
  reg [31:0] _RAND_4367;
  reg [31:0] _RAND_4368;
  reg [31:0] _RAND_4369;
  reg [31:0] _RAND_4370;
  reg [31:0] _RAND_4371;
  reg [31:0] _RAND_4372;
  reg [31:0] _RAND_4373;
  reg [31:0] _RAND_4374;
  reg [31:0] _RAND_4375;
  reg [31:0] _RAND_4376;
  reg [31:0] _RAND_4377;
  reg [31:0] _RAND_4378;
  reg [31:0] _RAND_4379;
  reg [31:0] _RAND_4380;
  reg [31:0] _RAND_4381;
  reg [31:0] _RAND_4382;
  reg [31:0] _RAND_4383;
  reg [31:0] _RAND_4384;
  reg [31:0] _RAND_4385;
  reg [31:0] _RAND_4386;
  reg [31:0] _RAND_4387;
  reg [31:0] _RAND_4388;
  reg [31:0] _RAND_4389;
  reg [31:0] _RAND_4390;
  reg [31:0] _RAND_4391;
  reg [31:0] _RAND_4392;
  reg [31:0] _RAND_4393;
  reg [31:0] _RAND_4394;
  reg [31:0] _RAND_4395;
  reg [31:0] _RAND_4396;
  reg [31:0] _RAND_4397;
  reg [31:0] _RAND_4398;
  reg [31:0] _RAND_4399;
  reg [31:0] _RAND_4400;
  reg [31:0] _RAND_4401;
  reg [31:0] _RAND_4402;
  reg [31:0] _RAND_4403;
  reg [31:0] _RAND_4404;
  reg [31:0] _RAND_4405;
  reg [31:0] _RAND_4406;
  reg [31:0] _RAND_4407;
  reg [31:0] _RAND_4408;
  reg [31:0] _RAND_4409;
  reg [31:0] _RAND_4410;
  reg [31:0] _RAND_4411;
  reg [31:0] _RAND_4412;
  reg [31:0] _RAND_4413;
  reg [31:0] _RAND_4414;
  reg [31:0] _RAND_4415;
  reg [31:0] _RAND_4416;
  reg [31:0] _RAND_4417;
  reg [31:0] _RAND_4418;
  reg [31:0] _RAND_4419;
  reg [31:0] _RAND_4420;
  reg [31:0] _RAND_4421;
  reg [31:0] _RAND_4422;
  reg [31:0] _RAND_4423;
  reg [31:0] _RAND_4424;
  reg [31:0] _RAND_4425;
  reg [31:0] _RAND_4426;
  reg [31:0] _RAND_4427;
  reg [31:0] _RAND_4428;
  reg [31:0] _RAND_4429;
  reg [31:0] _RAND_4430;
  reg [31:0] _RAND_4431;
  reg [31:0] _RAND_4432;
  reg [31:0] _RAND_4433;
  reg [31:0] _RAND_4434;
  reg [31:0] _RAND_4435;
  reg [31:0] _RAND_4436;
  reg [31:0] _RAND_4437;
  reg [31:0] _RAND_4438;
  reg [31:0] _RAND_4439;
  reg [31:0] _RAND_4440;
  reg [31:0] _RAND_4441;
  reg [31:0] _RAND_4442;
  reg [31:0] _RAND_4443;
  reg [31:0] _RAND_4444;
  reg [31:0] _RAND_4445;
  reg [31:0] _RAND_4446;
  reg [31:0] _RAND_4447;
  reg [31:0] _RAND_4448;
  reg [31:0] _RAND_4449;
  reg [31:0] _RAND_4450;
  reg [31:0] _RAND_4451;
  reg [31:0] _RAND_4452;
  reg [31:0] _RAND_4453;
  reg [31:0] _RAND_4454;
  reg [31:0] _RAND_4455;
  reg [31:0] _RAND_4456;
  reg [31:0] _RAND_4457;
  reg [31:0] _RAND_4458;
  reg [31:0] _RAND_4459;
  reg [31:0] _RAND_4460;
  reg [31:0] _RAND_4461;
  reg [31:0] _RAND_4462;
  reg [31:0] _RAND_4463;
  reg [31:0] _RAND_4464;
  reg [31:0] _RAND_4465;
  reg [31:0] _RAND_4466;
  reg [31:0] _RAND_4467;
  reg [31:0] _RAND_4468;
  reg [31:0] _RAND_4469;
  reg [31:0] _RAND_4470;
  reg [31:0] _RAND_4471;
  reg [31:0] _RAND_4472;
  reg [31:0] _RAND_4473;
  reg [31:0] _RAND_4474;
  reg [31:0] _RAND_4475;
  reg [31:0] _RAND_4476;
  reg [31:0] _RAND_4477;
  reg [31:0] _RAND_4478;
  reg [31:0] _RAND_4479;
  reg [31:0] _RAND_4480;
  reg [31:0] _RAND_4481;
  reg [31:0] _RAND_4482;
  reg [31:0] _RAND_4483;
  reg [31:0] _RAND_4484;
  reg [31:0] _RAND_4485;
  reg [31:0] _RAND_4486;
  reg [31:0] _RAND_4487;
  reg [31:0] _RAND_4488;
  reg [31:0] _RAND_4489;
  reg [31:0] _RAND_4490;
  reg [31:0] _RAND_4491;
  reg [31:0] _RAND_4492;
  reg [31:0] _RAND_4493;
  reg [31:0] _RAND_4494;
  reg [31:0] _RAND_4495;
  reg [31:0] _RAND_4496;
  reg [31:0] _RAND_4497;
  reg [31:0] _RAND_4498;
  reg [31:0] _RAND_4499;
  reg [31:0] _RAND_4500;
  reg [31:0] _RAND_4501;
  reg [31:0] _RAND_4502;
  reg [31:0] _RAND_4503;
  reg [31:0] _RAND_4504;
  reg [31:0] _RAND_4505;
  reg [31:0] _RAND_4506;
  reg [31:0] _RAND_4507;
  reg [31:0] _RAND_4508;
  reg [31:0] _RAND_4509;
  reg [31:0] _RAND_4510;
  reg [31:0] _RAND_4511;
  reg [31:0] _RAND_4512;
  reg [31:0] _RAND_4513;
  reg [31:0] _RAND_4514;
  reg [31:0] _RAND_4515;
  reg [31:0] _RAND_4516;
  reg [31:0] _RAND_4517;
  reg [31:0] _RAND_4518;
  reg [31:0] _RAND_4519;
  reg [31:0] _RAND_4520;
  reg [31:0] _RAND_4521;
  reg [31:0] _RAND_4522;
  reg [31:0] _RAND_4523;
  reg [31:0] _RAND_4524;
  reg [31:0] _RAND_4525;
  reg [31:0] _RAND_4526;
  reg [31:0] _RAND_4527;
  reg [31:0] _RAND_4528;
  reg [31:0] _RAND_4529;
  reg [31:0] _RAND_4530;
  reg [31:0] _RAND_4531;
  reg [31:0] _RAND_4532;
  reg [31:0] _RAND_4533;
  reg [31:0] _RAND_4534;
  reg [31:0] _RAND_4535;
  reg [31:0] _RAND_4536;
  reg [31:0] _RAND_4537;
  reg [31:0] _RAND_4538;
  reg [31:0] _RAND_4539;
  reg [31:0] _RAND_4540;
  reg [31:0] _RAND_4541;
  reg [31:0] _RAND_4542;
  reg [31:0] _RAND_4543;
  reg [31:0] _RAND_4544;
  reg [31:0] _RAND_4545;
  reg [31:0] _RAND_4546;
  reg [31:0] _RAND_4547;
  reg [31:0] _RAND_4548;
  reg [31:0] _RAND_4549;
  reg [31:0] _RAND_4550;
  reg [31:0] _RAND_4551;
  reg [31:0] _RAND_4552;
  reg [31:0] _RAND_4553;
  reg [31:0] _RAND_4554;
  reg [31:0] _RAND_4555;
  reg [31:0] _RAND_4556;
  reg [31:0] _RAND_4557;
  reg [31:0] _RAND_4558;
  reg [31:0] _RAND_4559;
  reg [31:0] _RAND_4560;
  reg [31:0] _RAND_4561;
  reg [31:0] _RAND_4562;
  reg [31:0] _RAND_4563;
  reg [31:0] _RAND_4564;
  reg [31:0] _RAND_4565;
  reg [31:0] _RAND_4566;
  reg [31:0] _RAND_4567;
  reg [31:0] _RAND_4568;
  reg [31:0] _RAND_4569;
  reg [31:0] _RAND_4570;
  reg [31:0] _RAND_4571;
  reg [31:0] _RAND_4572;
  reg [31:0] _RAND_4573;
  reg [31:0] _RAND_4574;
  reg [31:0] _RAND_4575;
  reg [31:0] _RAND_4576;
  reg [31:0] _RAND_4577;
  reg [31:0] _RAND_4578;
  reg [31:0] _RAND_4579;
  reg [31:0] _RAND_4580;
  reg [31:0] _RAND_4581;
  reg [31:0] _RAND_4582;
  reg [31:0] _RAND_4583;
  reg [31:0] _RAND_4584;
  reg [31:0] _RAND_4585;
  reg [31:0] _RAND_4586;
  reg [31:0] _RAND_4587;
  reg [31:0] _RAND_4588;
  reg [31:0] _RAND_4589;
  reg [31:0] _RAND_4590;
  reg [31:0] _RAND_4591;
  reg [31:0] _RAND_4592;
  reg [31:0] _RAND_4593;
  reg [31:0] _RAND_4594;
  reg [31:0] _RAND_4595;
  reg [31:0] _RAND_4596;
  reg [31:0] _RAND_4597;
  reg [31:0] _RAND_4598;
  reg [31:0] _RAND_4599;
  reg [31:0] _RAND_4600;
  reg [31:0] _RAND_4601;
  reg [31:0] _RAND_4602;
  reg [31:0] _RAND_4603;
  reg [31:0] _RAND_4604;
  reg [31:0] _RAND_4605;
  reg [31:0] _RAND_4606;
  reg [31:0] _RAND_4607;
  reg [31:0] _RAND_4608;
  reg [31:0] _RAND_4609;
  reg [31:0] _RAND_4610;
  reg [31:0] _RAND_4611;
  reg [31:0] _RAND_4612;
  reg [31:0] _RAND_4613;
  reg [31:0] _RAND_4614;
  reg [31:0] _RAND_4615;
  reg [31:0] _RAND_4616;
  reg [31:0] _RAND_4617;
  reg [31:0] _RAND_4618;
  reg [31:0] _RAND_4619;
  reg [31:0] _RAND_4620;
  reg [31:0] _RAND_4621;
  reg [31:0] _RAND_4622;
  reg [31:0] _RAND_4623;
  reg [31:0] _RAND_4624;
  reg [31:0] _RAND_4625;
  reg [31:0] _RAND_4626;
  reg [31:0] _RAND_4627;
  reg [31:0] _RAND_4628;
  reg [31:0] _RAND_4629;
  reg [31:0] _RAND_4630;
  reg [31:0] _RAND_4631;
  reg [31:0] _RAND_4632;
  reg [31:0] _RAND_4633;
  reg [31:0] _RAND_4634;
  reg [31:0] _RAND_4635;
  reg [31:0] _RAND_4636;
  reg [31:0] _RAND_4637;
  reg [31:0] _RAND_4638;
  reg [31:0] _RAND_4639;
  reg [31:0] _RAND_4640;
  reg [31:0] _RAND_4641;
  reg [31:0] _RAND_4642;
  reg [31:0] _RAND_4643;
  reg [31:0] _RAND_4644;
  reg [31:0] _RAND_4645;
  reg [31:0] _RAND_4646;
  reg [31:0] _RAND_4647;
  reg [31:0] _RAND_4648;
  reg [31:0] _RAND_4649;
  reg [31:0] _RAND_4650;
  reg [31:0] _RAND_4651;
  reg [31:0] _RAND_4652;
  reg [31:0] _RAND_4653;
  reg [31:0] _RAND_4654;
  reg [31:0] _RAND_4655;
  reg [31:0] _RAND_4656;
  reg [31:0] _RAND_4657;
  reg [31:0] _RAND_4658;
  reg [31:0] _RAND_4659;
  reg [31:0] _RAND_4660;
  reg [31:0] _RAND_4661;
  reg [31:0] _RAND_4662;
  reg [31:0] _RAND_4663;
  reg [31:0] _RAND_4664;
  reg [31:0] _RAND_4665;
  reg [31:0] _RAND_4666;
  reg [31:0] _RAND_4667;
  reg [31:0] _RAND_4668;
  reg [31:0] _RAND_4669;
  reg [31:0] _RAND_4670;
  reg [31:0] _RAND_4671;
  reg [31:0] _RAND_4672;
  reg [31:0] _RAND_4673;
  reg [31:0] _RAND_4674;
  reg [31:0] _RAND_4675;
  reg [31:0] _RAND_4676;
  reg [31:0] _RAND_4677;
  reg [31:0] _RAND_4678;
  reg [31:0] _RAND_4679;
  reg [31:0] _RAND_4680;
  reg [31:0] _RAND_4681;
  reg [31:0] _RAND_4682;
  reg [31:0] _RAND_4683;
  reg [31:0] _RAND_4684;
  reg [31:0] _RAND_4685;
  reg [31:0] _RAND_4686;
  reg [31:0] _RAND_4687;
  reg [31:0] _RAND_4688;
  reg [31:0] _RAND_4689;
  reg [31:0] _RAND_4690;
  reg [31:0] _RAND_4691;
  reg [31:0] _RAND_4692;
  reg [31:0] _RAND_4693;
  reg [31:0] _RAND_4694;
  reg [31:0] _RAND_4695;
  reg [31:0] _RAND_4696;
  reg [31:0] _RAND_4697;
  reg [31:0] _RAND_4698;
  reg [31:0] _RAND_4699;
  reg [31:0] _RAND_4700;
  reg [31:0] _RAND_4701;
  reg [31:0] _RAND_4702;
  reg [31:0] _RAND_4703;
  reg [31:0] _RAND_4704;
  reg [31:0] _RAND_4705;
  reg [31:0] _RAND_4706;
  reg [31:0] _RAND_4707;
  reg [31:0] _RAND_4708;
  reg [31:0] _RAND_4709;
  reg [31:0] _RAND_4710;
  reg [31:0] _RAND_4711;
  reg [31:0] _RAND_4712;
  reg [31:0] _RAND_4713;
  reg [31:0] _RAND_4714;
  reg [31:0] _RAND_4715;
  reg [31:0] _RAND_4716;
  reg [31:0] _RAND_4717;
  reg [31:0] _RAND_4718;
  reg [31:0] _RAND_4719;
  reg [31:0] _RAND_4720;
  reg [31:0] _RAND_4721;
  reg [31:0] _RAND_4722;
  reg [31:0] _RAND_4723;
  reg [31:0] _RAND_4724;
  reg [31:0] _RAND_4725;
  reg [31:0] _RAND_4726;
  reg [31:0] _RAND_4727;
  reg [31:0] _RAND_4728;
  reg [31:0] _RAND_4729;
  reg [31:0] _RAND_4730;
  reg [31:0] _RAND_4731;
  reg [31:0] _RAND_4732;
  reg [31:0] _RAND_4733;
  reg [31:0] _RAND_4734;
  reg [31:0] _RAND_4735;
  reg [31:0] _RAND_4736;
  reg [31:0] _RAND_4737;
  reg [31:0] _RAND_4738;
  reg [31:0] _RAND_4739;
  reg [31:0] _RAND_4740;
  reg [31:0] _RAND_4741;
  reg [31:0] _RAND_4742;
  reg [31:0] _RAND_4743;
  reg [31:0] _RAND_4744;
  reg [31:0] _RAND_4745;
  reg [31:0] _RAND_4746;
  reg [31:0] _RAND_4747;
  reg [31:0] _RAND_4748;
  reg [31:0] _RAND_4749;
  reg [31:0] _RAND_4750;
  reg [31:0] _RAND_4751;
  reg [31:0] _RAND_4752;
  reg [31:0] _RAND_4753;
  reg [31:0] _RAND_4754;
  reg [31:0] _RAND_4755;
  reg [31:0] _RAND_4756;
  reg [31:0] _RAND_4757;
  reg [31:0] _RAND_4758;
  reg [31:0] _RAND_4759;
  reg [31:0] _RAND_4760;
  reg [31:0] _RAND_4761;
  reg [31:0] _RAND_4762;
  reg [31:0] _RAND_4763;
  reg [31:0] _RAND_4764;
  reg [31:0] _RAND_4765;
  reg [31:0] _RAND_4766;
  reg [31:0] _RAND_4767;
  reg [31:0] _RAND_4768;
  reg [31:0] _RAND_4769;
  reg [31:0] _RAND_4770;
  reg [31:0] _RAND_4771;
  reg [31:0] _RAND_4772;
  reg [31:0] _RAND_4773;
  reg [31:0] _RAND_4774;
  reg [31:0] _RAND_4775;
  reg [31:0] _RAND_4776;
  reg [31:0] _RAND_4777;
  reg [31:0] _RAND_4778;
  reg [31:0] _RAND_4779;
  reg [31:0] _RAND_4780;
  reg [31:0] _RAND_4781;
  reg [31:0] _RAND_4782;
  reg [31:0] _RAND_4783;
  reg [31:0] _RAND_4784;
  reg [31:0] _RAND_4785;
  reg [31:0] _RAND_4786;
  reg [31:0] _RAND_4787;
  reg [31:0] _RAND_4788;
  reg [31:0] _RAND_4789;
  reg [31:0] _RAND_4790;
  reg [31:0] _RAND_4791;
  reg [31:0] _RAND_4792;
  reg [31:0] _RAND_4793;
  reg [31:0] _RAND_4794;
  reg [31:0] _RAND_4795;
  reg [31:0] _RAND_4796;
  reg [31:0] _RAND_4797;
  reg [31:0] _RAND_4798;
  reg [31:0] _RAND_4799;
  reg [31:0] _RAND_4800;
  reg [31:0] _RAND_4801;
  reg [31:0] _RAND_4802;
  reg [31:0] _RAND_4803;
  reg [31:0] _RAND_4804;
  reg [31:0] _RAND_4805;
  reg [31:0] _RAND_4806;
  reg [31:0] _RAND_4807;
  reg [31:0] _RAND_4808;
  reg [31:0] _RAND_4809;
  reg [31:0] _RAND_4810;
  reg [31:0] _RAND_4811;
  reg [31:0] _RAND_4812;
  reg [31:0] _RAND_4813;
  reg [31:0] _RAND_4814;
  reg [31:0] _RAND_4815;
  reg [31:0] _RAND_4816;
  reg [31:0] _RAND_4817;
  reg [31:0] _RAND_4818;
  reg [31:0] _RAND_4819;
  reg [31:0] _RAND_4820;
  reg [31:0] _RAND_4821;
  reg [31:0] _RAND_4822;
  reg [31:0] _RAND_4823;
  reg [31:0] _RAND_4824;
  reg [31:0] _RAND_4825;
  reg [31:0] _RAND_4826;
  reg [31:0] _RAND_4827;
  reg [31:0] _RAND_4828;
  reg [31:0] _RAND_4829;
  reg [31:0] _RAND_4830;
  reg [31:0] _RAND_4831;
  reg [31:0] _RAND_4832;
  reg [31:0] _RAND_4833;
  reg [31:0] _RAND_4834;
  reg [31:0] _RAND_4835;
  reg [31:0] _RAND_4836;
  reg [31:0] _RAND_4837;
  reg [31:0] _RAND_4838;
  reg [31:0] _RAND_4839;
  reg [31:0] _RAND_4840;
  reg [31:0] _RAND_4841;
  reg [31:0] _RAND_4842;
  reg [31:0] _RAND_4843;
  reg [31:0] _RAND_4844;
  reg [31:0] _RAND_4845;
  reg [31:0] _RAND_4846;
  reg [31:0] _RAND_4847;
  reg [31:0] _RAND_4848;
  reg [31:0] _RAND_4849;
  reg [31:0] _RAND_4850;
  reg [31:0] _RAND_4851;
  reg [31:0] _RAND_4852;
  reg [31:0] _RAND_4853;
  reg [31:0] _RAND_4854;
  reg [31:0] _RAND_4855;
  reg [31:0] _RAND_4856;
  reg [31:0] _RAND_4857;
  reg [31:0] _RAND_4858;
  reg [31:0] _RAND_4859;
  reg [31:0] _RAND_4860;
  reg [31:0] _RAND_4861;
  reg [31:0] _RAND_4862;
  reg [31:0] _RAND_4863;
  reg [31:0] _RAND_4864;
  reg [31:0] _RAND_4865;
  reg [31:0] _RAND_4866;
  reg [31:0] _RAND_4867;
  reg [31:0] _RAND_4868;
  reg [31:0] _RAND_4869;
  reg [31:0] _RAND_4870;
  reg [31:0] _RAND_4871;
  reg [31:0] _RAND_4872;
  reg [31:0] _RAND_4873;
  reg [31:0] _RAND_4874;
  reg [31:0] _RAND_4875;
  reg [31:0] _RAND_4876;
  reg [31:0] _RAND_4877;
  reg [31:0] _RAND_4878;
  reg [31:0] _RAND_4879;
  reg [31:0] _RAND_4880;
  reg [31:0] _RAND_4881;
  reg [31:0] _RAND_4882;
  reg [31:0] _RAND_4883;
  reg [31:0] _RAND_4884;
  reg [31:0] _RAND_4885;
  reg [31:0] _RAND_4886;
  reg [31:0] _RAND_4887;
  reg [31:0] _RAND_4888;
  reg [31:0] _RAND_4889;
  reg [31:0] _RAND_4890;
  reg [31:0] _RAND_4891;
  reg [31:0] _RAND_4892;
  reg [31:0] _RAND_4893;
  reg [31:0] _RAND_4894;
  reg [31:0] _RAND_4895;
  reg [31:0] _RAND_4896;
  reg [31:0] _RAND_4897;
  reg [31:0] _RAND_4898;
  reg [31:0] _RAND_4899;
  reg [31:0] _RAND_4900;
  reg [31:0] _RAND_4901;
  reg [31:0] _RAND_4902;
  reg [31:0] _RAND_4903;
  reg [31:0] _RAND_4904;
  reg [31:0] _RAND_4905;
  reg [31:0] _RAND_4906;
  reg [31:0] _RAND_4907;
  reg [31:0] _RAND_4908;
  reg [31:0] _RAND_4909;
  reg [31:0] _RAND_4910;
  reg [31:0] _RAND_4911;
  reg [31:0] _RAND_4912;
  reg [31:0] _RAND_4913;
  reg [31:0] _RAND_4914;
  reg [31:0] _RAND_4915;
  reg [31:0] _RAND_4916;
  reg [31:0] _RAND_4917;
  reg [31:0] _RAND_4918;
  reg [31:0] _RAND_4919;
  reg [31:0] _RAND_4920;
  reg [31:0] _RAND_4921;
  reg [31:0] _RAND_4922;
  reg [31:0] _RAND_4923;
  reg [31:0] _RAND_4924;
  reg [31:0] _RAND_4925;
  reg [31:0] _RAND_4926;
  reg [31:0] _RAND_4927;
  reg [31:0] _RAND_4928;
  reg [31:0] _RAND_4929;
  reg [31:0] _RAND_4930;
  reg [31:0] _RAND_4931;
  reg [31:0] _RAND_4932;
  reg [31:0] _RAND_4933;
  reg [31:0] _RAND_4934;
  reg [31:0] _RAND_4935;
  reg [31:0] _RAND_4936;
  reg [31:0] _RAND_4937;
  reg [31:0] _RAND_4938;
  reg [31:0] _RAND_4939;
  reg [31:0] _RAND_4940;
  reg [31:0] _RAND_4941;
  reg [31:0] _RAND_4942;
  reg [31:0] _RAND_4943;
  reg [31:0] _RAND_4944;
  reg [31:0] _RAND_4945;
  reg [31:0] _RAND_4946;
  reg [31:0] _RAND_4947;
  reg [31:0] _RAND_4948;
  reg [31:0] _RAND_4949;
  reg [31:0] _RAND_4950;
  reg [31:0] _RAND_4951;
  reg [31:0] _RAND_4952;
  reg [31:0] _RAND_4953;
  reg [31:0] _RAND_4954;
  reg [31:0] _RAND_4955;
  reg [31:0] _RAND_4956;
  reg [31:0] _RAND_4957;
  reg [31:0] _RAND_4958;
  reg [31:0] _RAND_4959;
  reg [31:0] _RAND_4960;
  reg [31:0] _RAND_4961;
  reg [31:0] _RAND_4962;
  reg [31:0] _RAND_4963;
  reg [31:0] _RAND_4964;
  reg [31:0] _RAND_4965;
  reg [31:0] _RAND_4966;
  reg [31:0] _RAND_4967;
  reg [31:0] _RAND_4968;
  reg [31:0] _RAND_4969;
  reg [31:0] _RAND_4970;
  reg [31:0] _RAND_4971;
  reg [31:0] _RAND_4972;
  reg [31:0] _RAND_4973;
  reg [31:0] _RAND_4974;
  reg [31:0] _RAND_4975;
  reg [31:0] _RAND_4976;
  reg [31:0] _RAND_4977;
  reg [31:0] _RAND_4978;
  reg [31:0] _RAND_4979;
  reg [31:0] _RAND_4980;
  reg [31:0] _RAND_4981;
  reg [31:0] _RAND_4982;
  reg [31:0] _RAND_4983;
  reg [31:0] _RAND_4984;
  reg [31:0] _RAND_4985;
  reg [31:0] _RAND_4986;
  reg [31:0] _RAND_4987;
  reg [31:0] _RAND_4988;
  reg [31:0] _RAND_4989;
  reg [31:0] _RAND_4990;
  reg [31:0] _RAND_4991;
  reg [31:0] _RAND_4992;
  reg [31:0] _RAND_4993;
  reg [31:0] _RAND_4994;
  reg [31:0] _RAND_4995;
  reg [31:0] _RAND_4996;
  reg [31:0] _RAND_4997;
  reg [31:0] _RAND_4998;
  reg [31:0] _RAND_4999;
  reg [31:0] _RAND_5000;
  reg [31:0] _RAND_5001;
  reg [31:0] _RAND_5002;
  reg [31:0] _RAND_5003;
  reg [31:0] _RAND_5004;
  reg [31:0] _RAND_5005;
  reg [31:0] _RAND_5006;
  reg [31:0] _RAND_5007;
  reg [31:0] _RAND_5008;
  reg [31:0] _RAND_5009;
  reg [31:0] _RAND_5010;
  reg [31:0] _RAND_5011;
  reg [31:0] _RAND_5012;
  reg [31:0] _RAND_5013;
  reg [31:0] _RAND_5014;
  reg [31:0] _RAND_5015;
  reg [31:0] _RAND_5016;
  reg [31:0] _RAND_5017;
  reg [31:0] _RAND_5018;
  reg [31:0] _RAND_5019;
  reg [31:0] _RAND_5020;
  reg [31:0] _RAND_5021;
  reg [31:0] _RAND_5022;
  reg [31:0] _RAND_5023;
  reg [31:0] _RAND_5024;
  reg [31:0] _RAND_5025;
  reg [31:0] _RAND_5026;
  reg [31:0] _RAND_5027;
  reg [31:0] _RAND_5028;
  reg [31:0] _RAND_5029;
  reg [31:0] _RAND_5030;
  reg [31:0] _RAND_5031;
  reg [31:0] _RAND_5032;
  reg [31:0] _RAND_5033;
  reg [31:0] _RAND_5034;
  reg [31:0] _RAND_5035;
  reg [31:0] _RAND_5036;
  reg [31:0] _RAND_5037;
  reg [31:0] _RAND_5038;
  reg [31:0] _RAND_5039;
  reg [31:0] _RAND_5040;
  reg [31:0] _RAND_5041;
  reg [31:0] _RAND_5042;
  reg [31:0] _RAND_5043;
  reg [31:0] _RAND_5044;
  reg [31:0] _RAND_5045;
  reg [31:0] _RAND_5046;
  reg [31:0] _RAND_5047;
  reg [31:0] _RAND_5048;
  reg [31:0] _RAND_5049;
  reg [31:0] _RAND_5050;
  reg [31:0] _RAND_5051;
  reg [31:0] _RAND_5052;
  reg [31:0] _RAND_5053;
  reg [31:0] _RAND_5054;
  reg [31:0] _RAND_5055;
  reg [31:0] _RAND_5056;
  reg [31:0] _RAND_5057;
  reg [31:0] _RAND_5058;
  reg [31:0] _RAND_5059;
  reg [31:0] _RAND_5060;
  reg [31:0] _RAND_5061;
  reg [31:0] _RAND_5062;
  reg [31:0] _RAND_5063;
  reg [31:0] _RAND_5064;
  reg [31:0] _RAND_5065;
  reg [31:0] _RAND_5066;
  reg [31:0] _RAND_5067;
  reg [31:0] _RAND_5068;
  reg [31:0] _RAND_5069;
  reg [31:0] _RAND_5070;
  reg [31:0] _RAND_5071;
  reg [31:0] _RAND_5072;
  reg [31:0] _RAND_5073;
  reg [31:0] _RAND_5074;
  reg [31:0] _RAND_5075;
  reg [31:0] _RAND_5076;
  reg [31:0] _RAND_5077;
  reg [31:0] _RAND_5078;
  reg [31:0] _RAND_5079;
  reg [31:0] _RAND_5080;
  reg [31:0] _RAND_5081;
  reg [31:0] _RAND_5082;
  reg [31:0] _RAND_5083;
  reg [31:0] _RAND_5084;
  reg [31:0] _RAND_5085;
  reg [31:0] _RAND_5086;
  reg [31:0] _RAND_5087;
  reg [31:0] _RAND_5088;
  reg [31:0] _RAND_5089;
  reg [31:0] _RAND_5090;
  reg [31:0] _RAND_5091;
  reg [31:0] _RAND_5092;
  reg [31:0] _RAND_5093;
  reg [31:0] _RAND_5094;
  reg [31:0] _RAND_5095;
  reg [31:0] _RAND_5096;
  reg [31:0] _RAND_5097;
  reg [31:0] _RAND_5098;
  reg [31:0] _RAND_5099;
  reg [31:0] _RAND_5100;
  reg [31:0] _RAND_5101;
  reg [31:0] _RAND_5102;
  reg [31:0] _RAND_5103;
  reg [31:0] _RAND_5104;
  reg [31:0] _RAND_5105;
  reg [31:0] _RAND_5106;
  reg [31:0] _RAND_5107;
  reg [31:0] _RAND_5108;
  reg [31:0] _RAND_5109;
  reg [31:0] _RAND_5110;
  reg [31:0] _RAND_5111;
  reg [31:0] _RAND_5112;
  reg [31:0] _RAND_5113;
  reg [31:0] _RAND_5114;
  reg [31:0] _RAND_5115;
  reg [31:0] _RAND_5116;
  reg [31:0] _RAND_5117;
  reg [31:0] _RAND_5118;
  reg [31:0] _RAND_5119;
  reg [31:0] _RAND_5120;
  reg [31:0] _RAND_5121;
  reg [31:0] _RAND_5122;
  reg [31:0] _RAND_5123;
  reg [31:0] _RAND_5124;
  reg [31:0] _RAND_5125;
  reg [31:0] _RAND_5126;
  reg [31:0] _RAND_5127;
  reg [31:0] _RAND_5128;
  reg [31:0] _RAND_5129;
  reg [31:0] _RAND_5130;
  reg [31:0] _RAND_5131;
  reg [31:0] _RAND_5132;
  reg [31:0] _RAND_5133;
  reg [31:0] _RAND_5134;
  reg [31:0] _RAND_5135;
  reg [31:0] _RAND_5136;
  reg [31:0] _RAND_5137;
  reg [31:0] _RAND_5138;
  reg [31:0] _RAND_5139;
  reg [31:0] _RAND_5140;
  reg [31:0] _RAND_5141;
  reg [31:0] _RAND_5142;
  reg [31:0] _RAND_5143;
  reg [31:0] _RAND_5144;
  reg [31:0] _RAND_5145;
  reg [31:0] _RAND_5146;
  reg [31:0] _RAND_5147;
  reg [31:0] _RAND_5148;
  reg [31:0] _RAND_5149;
  reg [31:0] _RAND_5150;
  reg [31:0] _RAND_5151;
  reg [31:0] _RAND_5152;
  reg [31:0] _RAND_5153;
  reg [31:0] _RAND_5154;
  reg [31:0] _RAND_5155;
  reg [31:0] _RAND_5156;
  reg [31:0] _RAND_5157;
  reg [31:0] _RAND_5158;
  reg [31:0] _RAND_5159;
  reg [31:0] _RAND_5160;
  reg [31:0] _RAND_5161;
  reg [31:0] _RAND_5162;
  reg [31:0] _RAND_5163;
  reg [31:0] _RAND_5164;
  reg [31:0] _RAND_5165;
  reg [31:0] _RAND_5166;
  reg [31:0] _RAND_5167;
  reg [31:0] _RAND_5168;
  reg [31:0] _RAND_5169;
  reg [31:0] _RAND_5170;
  reg [31:0] _RAND_5171;
  reg [31:0] _RAND_5172;
  reg [31:0] _RAND_5173;
  reg [31:0] _RAND_5174;
  reg [31:0] _RAND_5175;
  reg [31:0] _RAND_5176;
  reg [31:0] _RAND_5177;
  reg [31:0] _RAND_5178;
  reg [31:0] _RAND_5179;
  reg [31:0] _RAND_5180;
  reg [31:0] _RAND_5181;
  reg [31:0] _RAND_5182;
  reg [31:0] _RAND_5183;
  reg [31:0] _RAND_5184;
  reg [31:0] _RAND_5185;
  reg [31:0] _RAND_5186;
  reg [31:0] _RAND_5187;
  reg [31:0] _RAND_5188;
  reg [31:0] _RAND_5189;
  reg [31:0] _RAND_5190;
  reg [31:0] _RAND_5191;
  reg [31:0] _RAND_5192;
  reg [31:0] _RAND_5193;
  reg [31:0] _RAND_5194;
  reg [31:0] _RAND_5195;
  reg [31:0] _RAND_5196;
  reg [31:0] _RAND_5197;
  reg [31:0] _RAND_5198;
  reg [31:0] _RAND_5199;
  reg [31:0] _RAND_5200;
  reg [31:0] _RAND_5201;
  reg [31:0] _RAND_5202;
  reg [31:0] _RAND_5203;
  reg [31:0] _RAND_5204;
  reg [31:0] _RAND_5205;
  reg [31:0] _RAND_5206;
  reg [31:0] _RAND_5207;
  reg [31:0] _RAND_5208;
  reg [31:0] _RAND_5209;
  reg [31:0] _RAND_5210;
  reg [31:0] _RAND_5211;
  reg [31:0] _RAND_5212;
  reg [31:0] _RAND_5213;
  reg [31:0] _RAND_5214;
  reg [31:0] _RAND_5215;
  reg [31:0] _RAND_5216;
  reg [31:0] _RAND_5217;
  reg [31:0] _RAND_5218;
  reg [31:0] _RAND_5219;
  reg [31:0] _RAND_5220;
  reg [31:0] _RAND_5221;
  reg [31:0] _RAND_5222;
  reg [31:0] _RAND_5223;
  reg [31:0] _RAND_5224;
  reg [31:0] _RAND_5225;
  reg [31:0] _RAND_5226;
  reg [31:0] _RAND_5227;
  reg [31:0] _RAND_5228;
  reg [31:0] _RAND_5229;
  reg [31:0] _RAND_5230;
  reg [31:0] _RAND_5231;
  reg [31:0] _RAND_5232;
  reg [31:0] _RAND_5233;
  reg [31:0] _RAND_5234;
  reg [31:0] _RAND_5235;
  reg [31:0] _RAND_5236;
  reg [31:0] _RAND_5237;
  reg [31:0] _RAND_5238;
  reg [31:0] _RAND_5239;
  reg [31:0] _RAND_5240;
  reg [31:0] _RAND_5241;
  reg [31:0] _RAND_5242;
  reg [31:0] _RAND_5243;
  reg [31:0] _RAND_5244;
  reg [31:0] _RAND_5245;
  reg [31:0] _RAND_5246;
  reg [31:0] _RAND_5247;
  reg [31:0] _RAND_5248;
  reg [31:0] _RAND_5249;
  reg [31:0] _RAND_5250;
  reg [31:0] _RAND_5251;
  reg [31:0] _RAND_5252;
  reg [31:0] _RAND_5253;
  reg [31:0] _RAND_5254;
  reg [31:0] _RAND_5255;
  reg [31:0] _RAND_5256;
  reg [31:0] _RAND_5257;
  reg [31:0] _RAND_5258;
  reg [31:0] _RAND_5259;
  reg [31:0] _RAND_5260;
  reg [31:0] _RAND_5261;
  reg [31:0] _RAND_5262;
  reg [31:0] _RAND_5263;
  reg [31:0] _RAND_5264;
  reg [31:0] _RAND_5265;
  reg [31:0] _RAND_5266;
  reg [31:0] _RAND_5267;
  reg [31:0] _RAND_5268;
  reg [31:0] _RAND_5269;
  reg [31:0] _RAND_5270;
  reg [31:0] _RAND_5271;
  reg [31:0] _RAND_5272;
  reg [31:0] _RAND_5273;
  reg [31:0] _RAND_5274;
  reg [31:0] _RAND_5275;
  reg [31:0] _RAND_5276;
  reg [31:0] _RAND_5277;
  reg [31:0] _RAND_5278;
  reg [31:0] _RAND_5279;
  reg [31:0] _RAND_5280;
  reg [31:0] _RAND_5281;
  reg [31:0] _RAND_5282;
  reg [31:0] _RAND_5283;
  reg [31:0] _RAND_5284;
  reg [31:0] _RAND_5285;
  reg [31:0] _RAND_5286;
  reg [31:0] _RAND_5287;
  reg [31:0] _RAND_5288;
  reg [31:0] _RAND_5289;
  reg [31:0] _RAND_5290;
  reg [31:0] _RAND_5291;
  reg [31:0] _RAND_5292;
  reg [31:0] _RAND_5293;
  reg [31:0] _RAND_5294;
  reg [31:0] _RAND_5295;
  reg [31:0] _RAND_5296;
  reg [31:0] _RAND_5297;
  reg [31:0] _RAND_5298;
  reg [31:0] _RAND_5299;
  reg [31:0] _RAND_5300;
  reg [31:0] _RAND_5301;
  reg [31:0] _RAND_5302;
  reg [31:0] _RAND_5303;
  reg [31:0] _RAND_5304;
  reg [31:0] _RAND_5305;
  reg [31:0] _RAND_5306;
  reg [31:0] _RAND_5307;
  reg [31:0] _RAND_5308;
  reg [31:0] _RAND_5309;
  reg [31:0] _RAND_5310;
  reg [31:0] _RAND_5311;
  reg [31:0] _RAND_5312;
  reg [31:0] _RAND_5313;
  reg [31:0] _RAND_5314;
  reg [31:0] _RAND_5315;
  reg [31:0] _RAND_5316;
  reg [31:0] _RAND_5317;
  reg [31:0] _RAND_5318;
  reg [31:0] _RAND_5319;
  reg [31:0] _RAND_5320;
  reg [31:0] _RAND_5321;
  reg [31:0] _RAND_5322;
  reg [31:0] _RAND_5323;
  reg [31:0] _RAND_5324;
  reg [31:0] _RAND_5325;
  reg [31:0] _RAND_5326;
  reg [31:0] _RAND_5327;
  reg [31:0] _RAND_5328;
  reg [31:0] _RAND_5329;
  reg [31:0] _RAND_5330;
  reg [31:0] _RAND_5331;
  reg [31:0] _RAND_5332;
  reg [31:0] _RAND_5333;
  reg [31:0] _RAND_5334;
  reg [31:0] _RAND_5335;
  reg [31:0] _RAND_5336;
  reg [31:0] _RAND_5337;
  reg [31:0] _RAND_5338;
  reg [31:0] _RAND_5339;
  reg [31:0] _RAND_5340;
  reg [31:0] _RAND_5341;
  reg [31:0] _RAND_5342;
  reg [31:0] _RAND_5343;
  reg [31:0] _RAND_5344;
  reg [31:0] _RAND_5345;
  reg [31:0] _RAND_5346;
  reg [31:0] _RAND_5347;
  reg [31:0] _RAND_5348;
  reg [31:0] _RAND_5349;
  reg [31:0] _RAND_5350;
  reg [31:0] _RAND_5351;
  reg [31:0] _RAND_5352;
  reg [31:0] _RAND_5353;
  reg [31:0] _RAND_5354;
  reg [31:0] _RAND_5355;
  reg [31:0] _RAND_5356;
  reg [31:0] _RAND_5357;
  reg [31:0] _RAND_5358;
  reg [31:0] _RAND_5359;
  reg [31:0] _RAND_5360;
  reg [31:0] _RAND_5361;
  reg [31:0] _RAND_5362;
  reg [31:0] _RAND_5363;
  reg [31:0] _RAND_5364;
  reg [31:0] _RAND_5365;
  reg [31:0] _RAND_5366;
  reg [31:0] _RAND_5367;
  reg [31:0] _RAND_5368;
  reg [31:0] _RAND_5369;
  reg [31:0] _RAND_5370;
  reg [31:0] _RAND_5371;
  reg [31:0] _RAND_5372;
  reg [31:0] _RAND_5373;
  reg [31:0] _RAND_5374;
  reg [31:0] _RAND_5375;
  reg [31:0] _RAND_5376;
  reg [31:0] _RAND_5377;
  reg [31:0] _RAND_5378;
  reg [31:0] _RAND_5379;
  reg [31:0] _RAND_5380;
  reg [31:0] _RAND_5381;
  reg [31:0] _RAND_5382;
  reg [31:0] _RAND_5383;
  reg [31:0] _RAND_5384;
  reg [31:0] _RAND_5385;
  reg [31:0] _RAND_5386;
  reg [31:0] _RAND_5387;
  reg [31:0] _RAND_5388;
  reg [31:0] _RAND_5389;
  reg [31:0] _RAND_5390;
  reg [31:0] _RAND_5391;
  reg [31:0] _RAND_5392;
  reg [31:0] _RAND_5393;
  reg [31:0] _RAND_5394;
  reg [31:0] _RAND_5395;
  reg [31:0] _RAND_5396;
  reg [31:0] _RAND_5397;
  reg [31:0] _RAND_5398;
  reg [31:0] _RAND_5399;
  reg [31:0] _RAND_5400;
  reg [31:0] _RAND_5401;
  reg [31:0] _RAND_5402;
  reg [31:0] _RAND_5403;
  reg [31:0] _RAND_5404;
  reg [31:0] _RAND_5405;
  reg [31:0] _RAND_5406;
  reg [31:0] _RAND_5407;
  reg [31:0] _RAND_5408;
  reg [31:0] _RAND_5409;
  reg [31:0] _RAND_5410;
  reg [31:0] _RAND_5411;
  reg [31:0] _RAND_5412;
  reg [31:0] _RAND_5413;
  reg [31:0] _RAND_5414;
  reg [31:0] _RAND_5415;
  reg [31:0] _RAND_5416;
  reg [31:0] _RAND_5417;
  reg [31:0] _RAND_5418;
  reg [31:0] _RAND_5419;
  reg [31:0] _RAND_5420;
  reg [31:0] _RAND_5421;
  reg [31:0] _RAND_5422;
  reg [31:0] _RAND_5423;
  reg [31:0] _RAND_5424;
  reg [31:0] _RAND_5425;
  reg [31:0] _RAND_5426;
  reg [31:0] _RAND_5427;
  reg [31:0] _RAND_5428;
  reg [31:0] _RAND_5429;
  reg [31:0] _RAND_5430;
  reg [31:0] _RAND_5431;
  reg [31:0] _RAND_5432;
  reg [31:0] _RAND_5433;
  reg [31:0] _RAND_5434;
  reg [31:0] _RAND_5435;
  reg [31:0] _RAND_5436;
  reg [31:0] _RAND_5437;
  reg [31:0] _RAND_5438;
  reg [31:0] _RAND_5439;
  reg [31:0] _RAND_5440;
  reg [31:0] _RAND_5441;
  reg [31:0] _RAND_5442;
  reg [31:0] _RAND_5443;
  reg [31:0] _RAND_5444;
  reg [31:0] _RAND_5445;
  reg [31:0] _RAND_5446;
  reg [31:0] _RAND_5447;
  reg [31:0] _RAND_5448;
  reg [31:0] _RAND_5449;
  reg [31:0] _RAND_5450;
  reg [31:0] _RAND_5451;
  reg [31:0] _RAND_5452;
  reg [31:0] _RAND_5453;
  reg [31:0] _RAND_5454;
  reg [31:0] _RAND_5455;
  reg [31:0] _RAND_5456;
  reg [31:0] _RAND_5457;
  reg [31:0] _RAND_5458;
  reg [31:0] _RAND_5459;
  reg [31:0] _RAND_5460;
  reg [31:0] _RAND_5461;
  reg [31:0] _RAND_5462;
  reg [31:0] _RAND_5463;
  reg [31:0] _RAND_5464;
  reg [31:0] _RAND_5465;
  reg [31:0] _RAND_5466;
  reg [31:0] _RAND_5467;
  reg [31:0] _RAND_5468;
  reg [31:0] _RAND_5469;
  reg [31:0] _RAND_5470;
  reg [31:0] _RAND_5471;
  reg [31:0] _RAND_5472;
  reg [31:0] _RAND_5473;
  reg [31:0] _RAND_5474;
  reg [31:0] _RAND_5475;
  reg [31:0] _RAND_5476;
  reg [31:0] _RAND_5477;
  reg [31:0] _RAND_5478;
  reg [31:0] _RAND_5479;
  reg [31:0] _RAND_5480;
  reg [31:0] _RAND_5481;
  reg [31:0] _RAND_5482;
  reg [31:0] _RAND_5483;
  reg [31:0] _RAND_5484;
  reg [31:0] _RAND_5485;
  reg [31:0] _RAND_5486;
  reg [31:0] _RAND_5487;
  reg [31:0] _RAND_5488;
  reg [31:0] _RAND_5489;
  reg [31:0] _RAND_5490;
  reg [31:0] _RAND_5491;
  reg [31:0] _RAND_5492;
  reg [31:0] _RAND_5493;
  reg [31:0] _RAND_5494;
  reg [31:0] _RAND_5495;
  reg [31:0] _RAND_5496;
  reg [31:0] _RAND_5497;
  reg [31:0] _RAND_5498;
  reg [31:0] _RAND_5499;
  reg [31:0] _RAND_5500;
  reg [31:0] _RAND_5501;
  reg [31:0] _RAND_5502;
  reg [31:0] _RAND_5503;
  reg [31:0] _RAND_5504;
  reg [31:0] _RAND_5505;
  reg [31:0] _RAND_5506;
  reg [31:0] _RAND_5507;
  reg [31:0] _RAND_5508;
  reg [31:0] _RAND_5509;
  reg [31:0] _RAND_5510;
  reg [31:0] _RAND_5511;
  reg [31:0] _RAND_5512;
  reg [31:0] _RAND_5513;
  reg [31:0] _RAND_5514;
  reg [31:0] _RAND_5515;
  reg [31:0] _RAND_5516;
  reg [31:0] _RAND_5517;
  reg [31:0] _RAND_5518;
  reg [31:0] _RAND_5519;
  reg [31:0] _RAND_5520;
  reg [31:0] _RAND_5521;
  reg [31:0] _RAND_5522;
  reg [31:0] _RAND_5523;
  reg [31:0] _RAND_5524;
  reg [31:0] _RAND_5525;
  reg [31:0] _RAND_5526;
  reg [31:0] _RAND_5527;
  reg [31:0] _RAND_5528;
  reg [31:0] _RAND_5529;
  reg [31:0] _RAND_5530;
  reg [31:0] _RAND_5531;
  reg [31:0] _RAND_5532;
  reg [31:0] _RAND_5533;
  reg [31:0] _RAND_5534;
  reg [31:0] _RAND_5535;
  reg [31:0] _RAND_5536;
  reg [31:0] _RAND_5537;
  reg [31:0] _RAND_5538;
  reg [31:0] _RAND_5539;
  reg [31:0] _RAND_5540;
  reg [31:0] _RAND_5541;
  reg [31:0] _RAND_5542;
  reg [31:0] _RAND_5543;
  reg [31:0] _RAND_5544;
  reg [31:0] _RAND_5545;
  reg [31:0] _RAND_5546;
  reg [31:0] _RAND_5547;
  reg [31:0] _RAND_5548;
  reg [31:0] _RAND_5549;
  reg [31:0] _RAND_5550;
  reg [31:0] _RAND_5551;
  reg [31:0] _RAND_5552;
  reg [31:0] _RAND_5553;
  reg [31:0] _RAND_5554;
  reg [31:0] _RAND_5555;
  reg [31:0] _RAND_5556;
  reg [31:0] _RAND_5557;
  reg [31:0] _RAND_5558;
  reg [31:0] _RAND_5559;
  reg [31:0] _RAND_5560;
  reg [31:0] _RAND_5561;
  reg [31:0] _RAND_5562;
  reg [31:0] _RAND_5563;
  reg [31:0] _RAND_5564;
  reg [31:0] _RAND_5565;
  reg [31:0] _RAND_5566;
  reg [31:0] _RAND_5567;
  reg [31:0] _RAND_5568;
  reg [31:0] _RAND_5569;
  reg [31:0] _RAND_5570;
  reg [31:0] _RAND_5571;
  reg [31:0] _RAND_5572;
  reg [31:0] _RAND_5573;
  reg [31:0] _RAND_5574;
  reg [31:0] _RAND_5575;
  reg [31:0] _RAND_5576;
  reg [31:0] _RAND_5577;
  reg [31:0] _RAND_5578;
  reg [31:0] _RAND_5579;
  reg [31:0] _RAND_5580;
  reg [31:0] _RAND_5581;
  reg [31:0] _RAND_5582;
  reg [31:0] _RAND_5583;
  reg [31:0] _RAND_5584;
  reg [31:0] _RAND_5585;
  reg [31:0] _RAND_5586;
  reg [31:0] _RAND_5587;
  reg [31:0] _RAND_5588;
  reg [31:0] _RAND_5589;
  reg [31:0] _RAND_5590;
  reg [31:0] _RAND_5591;
  reg [31:0] _RAND_5592;
  reg [31:0] _RAND_5593;
  reg [31:0] _RAND_5594;
  reg [31:0] _RAND_5595;
  reg [31:0] _RAND_5596;
  reg [31:0] _RAND_5597;
  reg [31:0] _RAND_5598;
  reg [31:0] _RAND_5599;
  reg [31:0] _RAND_5600;
  reg [31:0] _RAND_5601;
  reg [31:0] _RAND_5602;
  reg [31:0] _RAND_5603;
  reg [31:0] _RAND_5604;
  reg [31:0] _RAND_5605;
  reg [31:0] _RAND_5606;
  reg [31:0] _RAND_5607;
  reg [31:0] _RAND_5608;
  reg [31:0] _RAND_5609;
  reg [31:0] _RAND_5610;
  reg [31:0] _RAND_5611;
  reg [31:0] _RAND_5612;
  reg [31:0] _RAND_5613;
  reg [31:0] _RAND_5614;
  reg [31:0] _RAND_5615;
  reg [31:0] _RAND_5616;
  reg [31:0] _RAND_5617;
  reg [31:0] _RAND_5618;
  reg [31:0] _RAND_5619;
  reg [31:0] _RAND_5620;
  reg [31:0] _RAND_5621;
  reg [31:0] _RAND_5622;
  reg [31:0] _RAND_5623;
  reg [31:0] _RAND_5624;
  reg [31:0] _RAND_5625;
  reg [31:0] _RAND_5626;
  reg [31:0] _RAND_5627;
  reg [31:0] _RAND_5628;
  reg [31:0] _RAND_5629;
  reg [31:0] _RAND_5630;
  reg [31:0] _RAND_5631;
  reg [31:0] _RAND_5632;
  reg [31:0] _RAND_5633;
  reg [31:0] _RAND_5634;
  reg [31:0] _RAND_5635;
  reg [31:0] _RAND_5636;
  reg [31:0] _RAND_5637;
  reg [31:0] _RAND_5638;
  reg [31:0] _RAND_5639;
  reg [31:0] _RAND_5640;
  reg [31:0] _RAND_5641;
  reg [31:0] _RAND_5642;
  reg [31:0] _RAND_5643;
  reg [31:0] _RAND_5644;
  reg [31:0] _RAND_5645;
  reg [31:0] _RAND_5646;
  reg [31:0] _RAND_5647;
  reg [31:0] _RAND_5648;
  reg [31:0] _RAND_5649;
  reg [31:0] _RAND_5650;
  reg [31:0] _RAND_5651;
  reg [31:0] _RAND_5652;
  reg [31:0] _RAND_5653;
  reg [31:0] _RAND_5654;
  reg [31:0] _RAND_5655;
  reg [31:0] _RAND_5656;
  reg [31:0] _RAND_5657;
  reg [31:0] _RAND_5658;
  reg [31:0] _RAND_5659;
  reg [31:0] _RAND_5660;
  reg [31:0] _RAND_5661;
  reg [31:0] _RAND_5662;
  reg [31:0] _RAND_5663;
  reg [31:0] _RAND_5664;
  reg [31:0] _RAND_5665;
  reg [31:0] _RAND_5666;
  reg [31:0] _RAND_5667;
  reg [31:0] _RAND_5668;
  reg [31:0] _RAND_5669;
  reg [31:0] _RAND_5670;
  reg [31:0] _RAND_5671;
  reg [31:0] _RAND_5672;
  reg [31:0] _RAND_5673;
  reg [31:0] _RAND_5674;
  reg [31:0] _RAND_5675;
  reg [31:0] _RAND_5676;
  reg [31:0] _RAND_5677;
  reg [31:0] _RAND_5678;
  reg [31:0] _RAND_5679;
  reg [31:0] _RAND_5680;
  reg [31:0] _RAND_5681;
  reg [31:0] _RAND_5682;
  reg [31:0] _RAND_5683;
  reg [31:0] _RAND_5684;
  reg [31:0] _RAND_5685;
  reg [31:0] _RAND_5686;
  reg [31:0] _RAND_5687;
  reg [31:0] _RAND_5688;
  reg [31:0] _RAND_5689;
  reg [31:0] _RAND_5690;
  reg [31:0] _RAND_5691;
  reg [31:0] _RAND_5692;
  reg [31:0] _RAND_5693;
  reg [31:0] _RAND_5694;
  reg [31:0] _RAND_5695;
  reg [31:0] _RAND_5696;
  reg [31:0] _RAND_5697;
  reg [31:0] _RAND_5698;
  reg [31:0] _RAND_5699;
  reg [31:0] _RAND_5700;
  reg [31:0] _RAND_5701;
  reg [31:0] _RAND_5702;
  reg [31:0] _RAND_5703;
  reg [31:0] _RAND_5704;
  reg [31:0] _RAND_5705;
  reg [31:0] _RAND_5706;
  reg [31:0] _RAND_5707;
  reg [31:0] _RAND_5708;
  reg [31:0] _RAND_5709;
  reg [31:0] _RAND_5710;
  reg [31:0] _RAND_5711;
  reg [31:0] _RAND_5712;
  reg [31:0] _RAND_5713;
  reg [31:0] _RAND_5714;
  reg [31:0] _RAND_5715;
  reg [31:0] _RAND_5716;
  reg [31:0] _RAND_5717;
  reg [31:0] _RAND_5718;
  reg [31:0] _RAND_5719;
  reg [31:0] _RAND_5720;
  reg [31:0] _RAND_5721;
  reg [31:0] _RAND_5722;
  reg [31:0] _RAND_5723;
  reg [31:0] _RAND_5724;
  reg [31:0] _RAND_5725;
  reg [31:0] _RAND_5726;
  reg [31:0] _RAND_5727;
  reg [31:0] _RAND_5728;
  reg [31:0] _RAND_5729;
  reg [31:0] _RAND_5730;
  reg [31:0] _RAND_5731;
  reg [31:0] _RAND_5732;
  reg [31:0] _RAND_5733;
  reg [31:0] _RAND_5734;
  reg [31:0] _RAND_5735;
  reg [31:0] _RAND_5736;
  reg [31:0] _RAND_5737;
  reg [31:0] _RAND_5738;
  reg [31:0] _RAND_5739;
  reg [31:0] _RAND_5740;
  reg [31:0] _RAND_5741;
  reg [31:0] _RAND_5742;
  reg [31:0] _RAND_5743;
  reg [31:0] _RAND_5744;
  reg [31:0] _RAND_5745;
  reg [31:0] _RAND_5746;
  reg [31:0] _RAND_5747;
  reg [31:0] _RAND_5748;
  reg [31:0] _RAND_5749;
  reg [31:0] _RAND_5750;
  reg [31:0] _RAND_5751;
  reg [31:0] _RAND_5752;
  reg [31:0] _RAND_5753;
  reg [31:0] _RAND_5754;
  reg [31:0] _RAND_5755;
  reg [31:0] _RAND_5756;
  reg [31:0] _RAND_5757;
  reg [31:0] _RAND_5758;
  reg [31:0] _RAND_5759;
  reg [31:0] _RAND_5760;
  reg [31:0] _RAND_5761;
  reg [31:0] _RAND_5762;
  reg [31:0] _RAND_5763;
  reg [31:0] _RAND_5764;
  reg [31:0] _RAND_5765;
  reg [31:0] _RAND_5766;
  reg [31:0] _RAND_5767;
  reg [31:0] _RAND_5768;
  reg [31:0] _RAND_5769;
  reg [31:0] _RAND_5770;
  reg [31:0] _RAND_5771;
  reg [31:0] _RAND_5772;
  reg [31:0] _RAND_5773;
  reg [31:0] _RAND_5774;
  reg [31:0] _RAND_5775;
  reg [31:0] _RAND_5776;
  reg [31:0] _RAND_5777;
  reg [31:0] _RAND_5778;
  reg [31:0] _RAND_5779;
  reg [31:0] _RAND_5780;
  reg [31:0] _RAND_5781;
  reg [31:0] _RAND_5782;
  reg [31:0] _RAND_5783;
  reg [31:0] _RAND_5784;
  reg [31:0] _RAND_5785;
  reg [31:0] _RAND_5786;
  reg [31:0] _RAND_5787;
  reg [31:0] _RAND_5788;
  reg [31:0] _RAND_5789;
  reg [31:0] _RAND_5790;
  reg [31:0] _RAND_5791;
  reg [31:0] _RAND_5792;
  reg [31:0] _RAND_5793;
  reg [31:0] _RAND_5794;
  reg [31:0] _RAND_5795;
  reg [31:0] _RAND_5796;
  reg [31:0] _RAND_5797;
  reg [31:0] _RAND_5798;
  reg [31:0] _RAND_5799;
  reg [31:0] _RAND_5800;
  reg [31:0] _RAND_5801;
  reg [31:0] _RAND_5802;
  reg [31:0] _RAND_5803;
  reg [31:0] _RAND_5804;
  reg [31:0] _RAND_5805;
  reg [31:0] _RAND_5806;
  reg [31:0] _RAND_5807;
  reg [31:0] _RAND_5808;
  reg [31:0] _RAND_5809;
  reg [31:0] _RAND_5810;
  reg [31:0] _RAND_5811;
  reg [31:0] _RAND_5812;
  reg [31:0] _RAND_5813;
  reg [31:0] _RAND_5814;
  reg [31:0] _RAND_5815;
  reg [31:0] _RAND_5816;
  reg [31:0] _RAND_5817;
  reg [31:0] _RAND_5818;
  reg [31:0] _RAND_5819;
  reg [31:0] _RAND_5820;
  reg [31:0] _RAND_5821;
  reg [31:0] _RAND_5822;
  reg [31:0] _RAND_5823;
  reg [31:0] _RAND_5824;
  reg [31:0] _RAND_5825;
  reg [31:0] _RAND_5826;
  reg [31:0] _RAND_5827;
  reg [31:0] _RAND_5828;
  reg [31:0] _RAND_5829;
  reg [31:0] _RAND_5830;
  reg [31:0] _RAND_5831;
  reg [31:0] _RAND_5832;
  reg [31:0] _RAND_5833;
  reg [31:0] _RAND_5834;
  reg [31:0] _RAND_5835;
  reg [31:0] _RAND_5836;
  reg [31:0] _RAND_5837;
  reg [31:0] _RAND_5838;
  reg [31:0] _RAND_5839;
  reg [31:0] _RAND_5840;
  reg [31:0] _RAND_5841;
  reg [31:0] _RAND_5842;
  reg [31:0] _RAND_5843;
  reg [31:0] _RAND_5844;
  reg [31:0] _RAND_5845;
  reg [31:0] _RAND_5846;
  reg [31:0] _RAND_5847;
  reg [31:0] _RAND_5848;
  reg [31:0] _RAND_5849;
  reg [31:0] _RAND_5850;
  reg [31:0] _RAND_5851;
  reg [31:0] _RAND_5852;
  reg [31:0] _RAND_5853;
  reg [31:0] _RAND_5854;
  reg [31:0] _RAND_5855;
  reg [31:0] _RAND_5856;
  reg [31:0] _RAND_5857;
  reg [31:0] _RAND_5858;
  reg [31:0] _RAND_5859;
  reg [31:0] _RAND_5860;
  reg [31:0] _RAND_5861;
  reg [31:0] _RAND_5862;
  reg [31:0] _RAND_5863;
  reg [31:0] _RAND_5864;
  reg [31:0] _RAND_5865;
  reg [31:0] _RAND_5866;
  reg [31:0] _RAND_5867;
  reg [31:0] _RAND_5868;
  reg [31:0] _RAND_5869;
  reg [31:0] _RAND_5870;
  reg [31:0] _RAND_5871;
  reg [31:0] _RAND_5872;
  reg [31:0] _RAND_5873;
  reg [31:0] _RAND_5874;
  reg [31:0] _RAND_5875;
  reg [31:0] _RAND_5876;
  reg [31:0] _RAND_5877;
  reg [31:0] _RAND_5878;
  reg [31:0] _RAND_5879;
  reg [31:0] _RAND_5880;
  reg [31:0] _RAND_5881;
  reg [31:0] _RAND_5882;
  reg [31:0] _RAND_5883;
  reg [31:0] _RAND_5884;
  reg [31:0] _RAND_5885;
  reg [31:0] _RAND_5886;
  reg [31:0] _RAND_5887;
  reg [31:0] _RAND_5888;
  reg [31:0] _RAND_5889;
  reg [31:0] _RAND_5890;
  reg [31:0] _RAND_5891;
  reg [31:0] _RAND_5892;
  reg [31:0] _RAND_5893;
  reg [31:0] _RAND_5894;
  reg [31:0] _RAND_5895;
  reg [31:0] _RAND_5896;
  reg [31:0] _RAND_5897;
  reg [31:0] _RAND_5898;
  reg [31:0] _RAND_5899;
  reg [31:0] _RAND_5900;
  reg [31:0] _RAND_5901;
  reg [31:0] _RAND_5902;
  reg [31:0] _RAND_5903;
  reg [31:0] _RAND_5904;
  reg [31:0] _RAND_5905;
  reg [31:0] _RAND_5906;
  reg [31:0] _RAND_5907;
  reg [31:0] _RAND_5908;
  reg [31:0] _RAND_5909;
  reg [31:0] _RAND_5910;
  reg [31:0] _RAND_5911;
  reg [31:0] _RAND_5912;
  reg [31:0] _RAND_5913;
  reg [31:0] _RAND_5914;
  reg [31:0] _RAND_5915;
  reg [31:0] _RAND_5916;
  reg [31:0] _RAND_5917;
  reg [31:0] _RAND_5918;
  reg [31:0] _RAND_5919;
  reg [31:0] _RAND_5920;
  reg [31:0] _RAND_5921;
  reg [31:0] _RAND_5922;
  reg [31:0] _RAND_5923;
  reg [31:0] _RAND_5924;
  reg [31:0] _RAND_5925;
  reg [31:0] _RAND_5926;
  reg [31:0] _RAND_5927;
  reg [31:0] _RAND_5928;
  reg [31:0] _RAND_5929;
  reg [31:0] _RAND_5930;
  reg [31:0] _RAND_5931;
  reg [31:0] _RAND_5932;
  reg [31:0] _RAND_5933;
  reg [31:0] _RAND_5934;
  reg [31:0] _RAND_5935;
  reg [31:0] _RAND_5936;
  reg [31:0] _RAND_5937;
  reg [31:0] _RAND_5938;
  reg [31:0] _RAND_5939;
  reg [31:0] _RAND_5940;
  reg [31:0] _RAND_5941;
  reg [31:0] _RAND_5942;
  reg [31:0] _RAND_5943;
  reg [31:0] _RAND_5944;
  reg [31:0] _RAND_5945;
  reg [31:0] _RAND_5946;
  reg [31:0] _RAND_5947;
  reg [31:0] _RAND_5948;
  reg [31:0] _RAND_5949;
  reg [31:0] _RAND_5950;
  reg [31:0] _RAND_5951;
  reg [31:0] _RAND_5952;
  reg [31:0] _RAND_5953;
  reg [31:0] _RAND_5954;
  reg [31:0] _RAND_5955;
  reg [31:0] _RAND_5956;
  reg [31:0] _RAND_5957;
  reg [31:0] _RAND_5958;
  reg [31:0] _RAND_5959;
  reg [31:0] _RAND_5960;
  reg [31:0] _RAND_5961;
  reg [31:0] _RAND_5962;
  reg [31:0] _RAND_5963;
  reg [31:0] _RAND_5964;
  reg [31:0] _RAND_5965;
  reg [31:0] _RAND_5966;
  reg [31:0] _RAND_5967;
  reg [31:0] _RAND_5968;
  reg [31:0] _RAND_5969;
  reg [31:0] _RAND_5970;
  reg [31:0] _RAND_5971;
  reg [31:0] _RAND_5972;
  reg [31:0] _RAND_5973;
  reg [31:0] _RAND_5974;
  reg [31:0] _RAND_5975;
  reg [31:0] _RAND_5976;
  reg [31:0] _RAND_5977;
  reg [31:0] _RAND_5978;
  reg [31:0] _RAND_5979;
  reg [31:0] _RAND_5980;
  reg [31:0] _RAND_5981;
  reg [31:0] _RAND_5982;
  reg [31:0] _RAND_5983;
  reg [31:0] _RAND_5984;
  reg [31:0] _RAND_5985;
  reg [31:0] _RAND_5986;
  reg [31:0] _RAND_5987;
  reg [31:0] _RAND_5988;
  reg [31:0] _RAND_5989;
  reg [31:0] _RAND_5990;
  reg [31:0] _RAND_5991;
  reg [31:0] _RAND_5992;
  reg [31:0] _RAND_5993;
  reg [31:0] _RAND_5994;
  reg [31:0] _RAND_5995;
  reg [31:0] _RAND_5996;
  reg [31:0] _RAND_5997;
  reg [31:0] _RAND_5998;
  reg [31:0] _RAND_5999;
  reg [31:0] _RAND_6000;
  reg [31:0] _RAND_6001;
  reg [31:0] _RAND_6002;
  reg [31:0] _RAND_6003;
  reg [31:0] _RAND_6004;
  reg [31:0] _RAND_6005;
  reg [31:0] _RAND_6006;
  reg [31:0] _RAND_6007;
  reg [31:0] _RAND_6008;
  reg [31:0] _RAND_6009;
  reg [31:0] _RAND_6010;
  reg [31:0] _RAND_6011;
  reg [31:0] _RAND_6012;
  reg [31:0] _RAND_6013;
  reg [31:0] _RAND_6014;
  reg [31:0] _RAND_6015;
  reg [31:0] _RAND_6016;
  reg [31:0] _RAND_6017;
  reg [31:0] _RAND_6018;
  reg [31:0] _RAND_6019;
  reg [31:0] _RAND_6020;
  reg [31:0] _RAND_6021;
  reg [31:0] _RAND_6022;
  reg [31:0] _RAND_6023;
  reg [31:0] _RAND_6024;
  reg [31:0] _RAND_6025;
  reg [31:0] _RAND_6026;
  reg [31:0] _RAND_6027;
  reg [31:0] _RAND_6028;
  reg [31:0] _RAND_6029;
  reg [31:0] _RAND_6030;
  reg [31:0] _RAND_6031;
  reg [31:0] _RAND_6032;
  reg [31:0] _RAND_6033;
  reg [31:0] _RAND_6034;
  reg [31:0] _RAND_6035;
  reg [31:0] _RAND_6036;
  reg [31:0] _RAND_6037;
  reg [31:0] _RAND_6038;
  reg [31:0] _RAND_6039;
  reg [31:0] _RAND_6040;
  reg [31:0] _RAND_6041;
  reg [31:0] _RAND_6042;
  reg [31:0] _RAND_6043;
  reg [31:0] _RAND_6044;
  reg [31:0] _RAND_6045;
  reg [31:0] _RAND_6046;
  reg [31:0] _RAND_6047;
  reg [31:0] _RAND_6048;
  reg [31:0] _RAND_6049;
  reg [31:0] _RAND_6050;
  reg [31:0] _RAND_6051;
  reg [31:0] _RAND_6052;
  reg [31:0] _RAND_6053;
  reg [31:0] _RAND_6054;
  reg [31:0] _RAND_6055;
  reg [31:0] _RAND_6056;
  reg [31:0] _RAND_6057;
  reg [31:0] _RAND_6058;
  reg [31:0] _RAND_6059;
  reg [31:0] _RAND_6060;
  reg [31:0] _RAND_6061;
  reg [31:0] _RAND_6062;
  reg [31:0] _RAND_6063;
  reg [31:0] _RAND_6064;
  reg [31:0] _RAND_6065;
  reg [31:0] _RAND_6066;
  reg [31:0] _RAND_6067;
  reg [31:0] _RAND_6068;
  reg [31:0] _RAND_6069;
  reg [31:0] _RAND_6070;
  reg [31:0] _RAND_6071;
  reg [31:0] _RAND_6072;
  reg [31:0] _RAND_6073;
  reg [31:0] _RAND_6074;
  reg [31:0] _RAND_6075;
  reg [31:0] _RAND_6076;
  reg [31:0] _RAND_6077;
  reg [31:0] _RAND_6078;
  reg [31:0] _RAND_6079;
  reg [31:0] _RAND_6080;
  reg [31:0] _RAND_6081;
  reg [31:0] _RAND_6082;
  reg [31:0] _RAND_6083;
  reg [31:0] _RAND_6084;
  reg [31:0] _RAND_6085;
  reg [31:0] _RAND_6086;
  reg [31:0] _RAND_6087;
  reg [31:0] _RAND_6088;
  reg [31:0] _RAND_6089;
  reg [31:0] _RAND_6090;
  reg [31:0] _RAND_6091;
  reg [31:0] _RAND_6092;
  reg [31:0] _RAND_6093;
  reg [31:0] _RAND_6094;
  reg [31:0] _RAND_6095;
  reg [31:0] _RAND_6096;
  reg [31:0] _RAND_6097;
  reg [31:0] _RAND_6098;
  reg [31:0] _RAND_6099;
  reg [31:0] _RAND_6100;
  reg [31:0] _RAND_6101;
  reg [31:0] _RAND_6102;
  reg [31:0] _RAND_6103;
  reg [31:0] _RAND_6104;
  reg [31:0] _RAND_6105;
  reg [31:0] _RAND_6106;
  reg [31:0] _RAND_6107;
  reg [31:0] _RAND_6108;
  reg [31:0] _RAND_6109;
  reg [31:0] _RAND_6110;
  reg [31:0] _RAND_6111;
  reg [31:0] _RAND_6112;
  reg [31:0] _RAND_6113;
  reg [31:0] _RAND_6114;
  reg [31:0] _RAND_6115;
  reg [31:0] _RAND_6116;
  reg [31:0] _RAND_6117;
  reg [31:0] _RAND_6118;
  reg [31:0] _RAND_6119;
  reg [31:0] _RAND_6120;
  reg [31:0] _RAND_6121;
  reg [31:0] _RAND_6122;
  reg [31:0] _RAND_6123;
  reg [31:0] _RAND_6124;
  reg [31:0] _RAND_6125;
  reg [31:0] _RAND_6126;
  reg [31:0] _RAND_6127;
  reg [31:0] _RAND_6128;
  reg [31:0] _RAND_6129;
  reg [31:0] _RAND_6130;
  reg [31:0] _RAND_6131;
  reg [31:0] _RAND_6132;
  reg [31:0] _RAND_6133;
  reg [31:0] _RAND_6134;
  reg [31:0] _RAND_6135;
  reg [31:0] _RAND_6136;
  reg [31:0] _RAND_6137;
  reg [31:0] _RAND_6138;
  reg [31:0] _RAND_6139;
  reg [31:0] _RAND_6140;
  reg [31:0] _RAND_6141;
  reg [31:0] _RAND_6142;
  reg [31:0] _RAND_6143;
  reg [31:0] _RAND_6144;
  reg [31:0] _RAND_6145;
  reg [31:0] _RAND_6146;
  reg [31:0] _RAND_6147;
  reg [31:0] _RAND_6148;
  reg [31:0] _RAND_6149;
  reg [31:0] _RAND_6150;
  reg [31:0] _RAND_6151;
  reg [31:0] _RAND_6152;
  reg [31:0] _RAND_6153;
  reg [31:0] _RAND_6154;
  reg [31:0] _RAND_6155;
  reg [31:0] _RAND_6156;
  reg [31:0] _RAND_6157;
  reg [31:0] _RAND_6158;
  reg [31:0] _RAND_6159;
  reg [31:0] _RAND_6160;
  reg [31:0] _RAND_6161;
  reg [31:0] _RAND_6162;
  reg [31:0] _RAND_6163;
  reg [31:0] _RAND_6164;
  reg [31:0] _RAND_6165;
  reg [31:0] _RAND_6166;
  reg [31:0] _RAND_6167;
  reg [31:0] _RAND_6168;
  reg [31:0] _RAND_6169;
  reg [31:0] _RAND_6170;
  reg [31:0] _RAND_6171;
  reg [31:0] _RAND_6172;
  reg [31:0] _RAND_6173;
  reg [31:0] _RAND_6174;
  reg [31:0] _RAND_6175;
  reg [31:0] _RAND_6176;
  reg [31:0] _RAND_6177;
  reg [31:0] _RAND_6178;
  reg [31:0] _RAND_6179;
  reg [31:0] _RAND_6180;
  reg [31:0] _RAND_6181;
  reg [31:0] _RAND_6182;
  reg [31:0] _RAND_6183;
  reg [31:0] _RAND_6184;
  reg [31:0] _RAND_6185;
  reg [31:0] _RAND_6186;
  reg [31:0] _RAND_6187;
  reg [31:0] _RAND_6188;
  reg [31:0] _RAND_6189;
  reg [31:0] _RAND_6190;
  reg [31:0] _RAND_6191;
  reg [31:0] _RAND_6192;
  reg [31:0] _RAND_6193;
  reg [31:0] _RAND_6194;
  reg [31:0] _RAND_6195;
  reg [31:0] _RAND_6196;
  reg [31:0] _RAND_6197;
  reg [31:0] _RAND_6198;
  reg [31:0] _RAND_6199;
  reg [31:0] _RAND_6200;
  reg [31:0] _RAND_6201;
  reg [31:0] _RAND_6202;
  reg [31:0] _RAND_6203;
  reg [31:0] _RAND_6204;
  reg [31:0] _RAND_6205;
  reg [31:0] _RAND_6206;
  reg [31:0] _RAND_6207;
  reg [31:0] _RAND_6208;
  reg [31:0] _RAND_6209;
  reg [31:0] _RAND_6210;
  reg [31:0] _RAND_6211;
  reg [31:0] _RAND_6212;
  reg [31:0] _RAND_6213;
  reg [31:0] _RAND_6214;
  reg [31:0] _RAND_6215;
  reg [31:0] _RAND_6216;
  reg [31:0] _RAND_6217;
  reg [31:0] _RAND_6218;
  reg [31:0] _RAND_6219;
  reg [31:0] _RAND_6220;
  reg [31:0] _RAND_6221;
  reg [31:0] _RAND_6222;
  reg [31:0] _RAND_6223;
  reg [31:0] _RAND_6224;
  reg [31:0] _RAND_6225;
  reg [31:0] _RAND_6226;
  reg [31:0] _RAND_6227;
  reg [31:0] _RAND_6228;
  reg [31:0] _RAND_6229;
  reg [31:0] _RAND_6230;
  reg [31:0] _RAND_6231;
  reg [31:0] _RAND_6232;
  reg [31:0] _RAND_6233;
  reg [31:0] _RAND_6234;
  reg [31:0] _RAND_6235;
  reg [31:0] _RAND_6236;
  reg [31:0] _RAND_6237;
  reg [31:0] _RAND_6238;
  reg [31:0] _RAND_6239;
  reg [31:0] _RAND_6240;
  reg [31:0] _RAND_6241;
  reg [31:0] _RAND_6242;
  reg [31:0] _RAND_6243;
  reg [31:0] _RAND_6244;
  reg [31:0] _RAND_6245;
  reg [31:0] _RAND_6246;
  reg [31:0] _RAND_6247;
  reg [31:0] _RAND_6248;
  reg [31:0] _RAND_6249;
  reg [31:0] _RAND_6250;
  reg [31:0] _RAND_6251;
  reg [31:0] _RAND_6252;
  reg [31:0] _RAND_6253;
  reg [31:0] _RAND_6254;
  reg [31:0] _RAND_6255;
  reg [31:0] _RAND_6256;
  reg [31:0] _RAND_6257;
  reg [31:0] _RAND_6258;
  reg [31:0] _RAND_6259;
  reg [31:0] _RAND_6260;
  reg [31:0] _RAND_6261;
  reg [31:0] _RAND_6262;
  reg [31:0] _RAND_6263;
  reg [31:0] _RAND_6264;
  reg [31:0] _RAND_6265;
  reg [31:0] _RAND_6266;
  reg [31:0] _RAND_6267;
  reg [31:0] _RAND_6268;
  reg [31:0] _RAND_6269;
  reg [31:0] _RAND_6270;
  reg [31:0] _RAND_6271;
  reg [31:0] _RAND_6272;
  reg [31:0] _RAND_6273;
  reg [31:0] _RAND_6274;
  reg [31:0] _RAND_6275;
  reg [31:0] _RAND_6276;
  reg [31:0] _RAND_6277;
  reg [31:0] _RAND_6278;
  reg [31:0] _RAND_6279;
  reg [31:0] _RAND_6280;
  reg [31:0] _RAND_6281;
  reg [31:0] _RAND_6282;
  reg [31:0] _RAND_6283;
  reg [31:0] _RAND_6284;
  reg [31:0] _RAND_6285;
  reg [31:0] _RAND_6286;
  reg [31:0] _RAND_6287;
  reg [31:0] _RAND_6288;
  reg [31:0] _RAND_6289;
  reg [31:0] _RAND_6290;
  reg [31:0] _RAND_6291;
  reg [31:0] _RAND_6292;
  reg [31:0] _RAND_6293;
  reg [31:0] _RAND_6294;
  reg [31:0] _RAND_6295;
  reg [31:0] _RAND_6296;
  reg [31:0] _RAND_6297;
  reg [31:0] _RAND_6298;
  reg [31:0] _RAND_6299;
  reg [31:0] _RAND_6300;
  reg [31:0] _RAND_6301;
  reg [31:0] _RAND_6302;
  reg [31:0] _RAND_6303;
  reg [31:0] _RAND_6304;
  reg [31:0] _RAND_6305;
  reg [31:0] _RAND_6306;
  reg [31:0] _RAND_6307;
  reg [31:0] _RAND_6308;
  reg [31:0] _RAND_6309;
  reg [31:0] _RAND_6310;
  reg [31:0] _RAND_6311;
  reg [31:0] _RAND_6312;
  reg [31:0] _RAND_6313;
  reg [31:0] _RAND_6314;
  reg [31:0] _RAND_6315;
  reg [31:0] _RAND_6316;
  reg [31:0] _RAND_6317;
  reg [31:0] _RAND_6318;
  reg [31:0] _RAND_6319;
  reg [31:0] _RAND_6320;
  reg [31:0] _RAND_6321;
  reg [31:0] _RAND_6322;
  reg [31:0] _RAND_6323;
  reg [31:0] _RAND_6324;
  reg [31:0] _RAND_6325;
  reg [31:0] _RAND_6326;
  reg [31:0] _RAND_6327;
  reg [31:0] _RAND_6328;
  reg [31:0] _RAND_6329;
  reg [31:0] _RAND_6330;
  reg [31:0] _RAND_6331;
  reg [31:0] _RAND_6332;
  reg [31:0] _RAND_6333;
  reg [31:0] _RAND_6334;
  reg [31:0] _RAND_6335;
  reg [31:0] _RAND_6336;
  reg [31:0] _RAND_6337;
  reg [31:0] _RAND_6338;
  reg [31:0] _RAND_6339;
  reg [31:0] _RAND_6340;
  reg [31:0] _RAND_6341;
  reg [31:0] _RAND_6342;
  reg [31:0] _RAND_6343;
  reg [31:0] _RAND_6344;
  reg [31:0] _RAND_6345;
  reg [31:0] _RAND_6346;
  reg [31:0] _RAND_6347;
  reg [31:0] _RAND_6348;
  reg [31:0] _RAND_6349;
  reg [31:0] _RAND_6350;
  reg [31:0] _RAND_6351;
  reg [31:0] _RAND_6352;
  reg [31:0] _RAND_6353;
  reg [31:0] _RAND_6354;
  reg [31:0] _RAND_6355;
  reg [31:0] _RAND_6356;
  reg [31:0] _RAND_6357;
  reg [31:0] _RAND_6358;
  reg [31:0] _RAND_6359;
  reg [31:0] _RAND_6360;
  reg [31:0] _RAND_6361;
  reg [31:0] _RAND_6362;
  reg [31:0] _RAND_6363;
  reg [31:0] _RAND_6364;
  reg [31:0] _RAND_6365;
  reg [31:0] _RAND_6366;
  reg [31:0] _RAND_6367;
  reg [31:0] _RAND_6368;
  reg [31:0] _RAND_6369;
  reg [31:0] _RAND_6370;
  reg [31:0] _RAND_6371;
  reg [31:0] _RAND_6372;
  reg [31:0] _RAND_6373;
  reg [31:0] _RAND_6374;
  reg [31:0] _RAND_6375;
  reg [31:0] _RAND_6376;
  reg [31:0] _RAND_6377;
  reg [31:0] _RAND_6378;
  reg [31:0] _RAND_6379;
  reg [31:0] _RAND_6380;
  reg [31:0] _RAND_6381;
  reg [31:0] _RAND_6382;
  reg [31:0] _RAND_6383;
  reg [31:0] _RAND_6384;
  reg [31:0] _RAND_6385;
  reg [31:0] _RAND_6386;
  reg [31:0] _RAND_6387;
  reg [31:0] _RAND_6388;
  reg [31:0] _RAND_6389;
  reg [31:0] _RAND_6390;
  reg [31:0] _RAND_6391;
  reg [31:0] _RAND_6392;
  reg [31:0] _RAND_6393;
  reg [31:0] _RAND_6394;
  reg [31:0] _RAND_6395;
  reg [31:0] _RAND_6396;
  reg [31:0] _RAND_6397;
  reg [31:0] _RAND_6398;
  reg [31:0] _RAND_6399;
  reg [31:0] _RAND_6400;
  reg [31:0] _RAND_6401;
  reg [31:0] _RAND_6402;
  reg [31:0] _RAND_6403;
  reg [31:0] _RAND_6404;
  reg [31:0] _RAND_6405;
  reg [31:0] _RAND_6406;
  reg [31:0] _RAND_6407;
  reg [31:0] _RAND_6408;
  reg [31:0] _RAND_6409;
  reg [31:0] _RAND_6410;
  reg [31:0] _RAND_6411;
  reg [31:0] _RAND_6412;
  reg [31:0] _RAND_6413;
  reg [31:0] _RAND_6414;
  reg [31:0] _RAND_6415;
  reg [31:0] _RAND_6416;
  reg [31:0] _RAND_6417;
  reg [31:0] _RAND_6418;
  reg [31:0] _RAND_6419;
  reg [31:0] _RAND_6420;
  reg [31:0] _RAND_6421;
  reg [31:0] _RAND_6422;
  reg [31:0] _RAND_6423;
  reg [31:0] _RAND_6424;
  reg [31:0] _RAND_6425;
  reg [31:0] _RAND_6426;
  reg [31:0] _RAND_6427;
  reg [31:0] _RAND_6428;
  reg [31:0] _RAND_6429;
  reg [31:0] _RAND_6430;
  reg [31:0] _RAND_6431;
`endif // RANDOMIZE_REG_INIT
  wire [7:0] MulAdd_io_b_0; // @[ChiselImProc.scala 206:29]
  wire [7:0] MulAdd_io_b_1; // @[ChiselImProc.scala 206:29]
  wire [7:0] MulAdd_io_b_2; // @[ChiselImProc.scala 206:29]
  wire [7:0] MulAdd_io_b_3; // @[ChiselImProc.scala 206:29]
  wire [7:0] MulAdd_io_b_4; // @[ChiselImProc.scala 206:29]
  wire [7:0] MulAdd_io_b_5; // @[ChiselImProc.scala 206:29]
  wire [7:0] MulAdd_io_b_6; // @[ChiselImProc.scala 206:29]
  wire [7:0] MulAdd_io_b_7; // @[ChiselImProc.scala 206:29]
  wire [7:0] MulAdd_io_b_8; // @[ChiselImProc.scala 206:29]
  wire [7:0] MulAdd_io_b_9; // @[ChiselImProc.scala 206:29]
  wire [7:0] MulAdd_io_b_10; // @[ChiselImProc.scala 206:29]
  wire [7:0] MulAdd_io_b_11; // @[ChiselImProc.scala 206:29]
  wire [7:0] MulAdd_io_b_12; // @[ChiselImProc.scala 206:29]
  wire [7:0] MulAdd_io_b_13; // @[ChiselImProc.scala 206:29]
  wire [7:0] MulAdd_io_b_14; // @[ChiselImProc.scala 206:29]
  wire [7:0] MulAdd_io_b_15; // @[ChiselImProc.scala 206:29]
  wire [7:0] MulAdd_io_b_16; // @[ChiselImProc.scala 206:29]
  wire [7:0] MulAdd_io_b_17; // @[ChiselImProc.scala 206:29]
  wire [7:0] MulAdd_io_b_18; // @[ChiselImProc.scala 206:29]
  wire [7:0] MulAdd_io_b_19; // @[ChiselImProc.scala 206:29]
  wire [7:0] MulAdd_io_b_20; // @[ChiselImProc.scala 206:29]
  wire [7:0] MulAdd_io_b_21; // @[ChiselImProc.scala 206:29]
  wire [7:0] MulAdd_io_b_22; // @[ChiselImProc.scala 206:29]
  wire [7:0] MulAdd_io_b_23; // @[ChiselImProc.scala 206:29]
  wire [7:0] MulAdd_io_b_24; // @[ChiselImProc.scala 206:29]
  wire [15:0] MulAdd_io_output; // @[ChiselImProc.scala 206:29]
  reg [1:0] stateReg; // @[ChiselImProc.scala 56:28]
  reg [7:0] dataReg; // @[ChiselImProc.scala 58:23]
  reg [7:0] shadowReg; // @[ChiselImProc.scala 60:25]
  reg  userReg; // @[ChiselImProc.scala 61:23]
  reg  shadowUserReg; // @[ChiselImProc.scala 62:29]
  reg  lastReg; // @[ChiselImProc.scala 63:23]
  reg  shadowLastReg; // @[ChiselImProc.scala 64:29]
  wire  _T = 2'h0 == stateReg; // @[Conditional.scala 37:30]
  wire  _T_1 = 2'h1 == stateReg; // @[Conditional.scala 37:30]
  wire  _T_2 = ~io_enq_valid; // @[ChiselImProc.scala 78:39]
  wire  _T_3 = io_deq_ready & _T_2; // @[ChiselImProc.scala 78:36]
  wire  _T_4 = io_deq_ready & io_enq_valid; // @[ChiselImProc.scala 81:42]
  wire  _T_5 = ~io_deq_ready; // @[ChiselImProc.scala 86:29]
  wire  _T_6 = _T_5 & io_enq_valid; // @[ChiselImProc.scala 86:43]
  wire  _T_7 = 2'h2 == stateReg; // @[Conditional.scala 37:30]
  wire  _T_8 = 2'h3 == stateReg; // @[Conditional.scala 37:30]
  wire  _T_9 = stateReg == 2'h0; // @[ChiselImProc.scala 110:35]
  wire  _T_10 = stateReg == 2'h1; // @[ChiselImProc.scala 110:57]
  wire  _T_11 = _T_9 | _T_10; // @[ChiselImProc.scala 110:45]
  wire  _T_12 = stateReg == 2'h3; // @[ChiselImProc.scala 110:77]
  wire  _T_15 = stateReg == 2'h2; // @[ChiselImProc.scala 111:55]
  wire  _T_16 = _T_10 | _T_15; // @[ChiselImProc.scala 111:43]
  reg [7:0] lineBuffer_0; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_6; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_7; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_8; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_9; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_10; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_11; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_12; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_13; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_14; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_15; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_16; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_17; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_18; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_19; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_20; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_21; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_22; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_23; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_24; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_25; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_26; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_27; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_28; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_29; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_30; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_31; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_32; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_33; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_34; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_35; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_36; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_37; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_38; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_39; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_40; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_41; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_42; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_43; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_44; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_45; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_46; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_47; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_48; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_49; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_50; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_51; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_52; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_53; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_54; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_55; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_56; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_57; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_58; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_59; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_60; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_61; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_62; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_63; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_64; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_65; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_66; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_67; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_68; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_69; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_70; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_71; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_72; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_73; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_74; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_75; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_76; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_77; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_78; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_79; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_80; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_81; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_82; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_83; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_84; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_85; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_86; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_87; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_88; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_89; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_90; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_91; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_92; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_93; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_94; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_95; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_96; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_97; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_98; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_99; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_100; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_101; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_102; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_103; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_104; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_105; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_106; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_107; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_108; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_109; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_110; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_111; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_112; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_113; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_114; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_115; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_116; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_117; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_118; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_119; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_120; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_121; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_122; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_123; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_124; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_125; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_126; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_127; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_128; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_129; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_130; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_131; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_132; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_133; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_134; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_135; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_136; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_137; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_138; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_139; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_140; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_141; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_142; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_143; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_144; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_145; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_146; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_147; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_148; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_149; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_150; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_151; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_152; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_153; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_154; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_155; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_156; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_157; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_158; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_159; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_160; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_161; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_162; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_163; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_164; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_165; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_166; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_167; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_168; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_169; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_170; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_171; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_172; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_173; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_174; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_175; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_176; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_177; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_178; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_179; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_180; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_181; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_182; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_183; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_184; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_185; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_186; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_187; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_188; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_189; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_190; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_191; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_192; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_193; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_194; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_195; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_196; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_197; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_198; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_199; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_200; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_201; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_202; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_203; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_204; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_205; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_206; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_207; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_208; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_209; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_210; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_211; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_212; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_213; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_214; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_215; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_216; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_217; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_218; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_219; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_220; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_221; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_222; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_223; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_224; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_225; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_226; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_227; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_228; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_229; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_230; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_231; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_232; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_233; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_234; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_235; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_236; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_237; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_238; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_239; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_240; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_241; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_242; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_243; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_244; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_245; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_246; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_247; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_248; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_249; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_250; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_251; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_252; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_253; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_254; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_255; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_256; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_257; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_258; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_259; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_260; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_261; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_262; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_263; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_264; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_265; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_266; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_267; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_268; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_269; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_270; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_271; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_272; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_273; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_274; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_275; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_276; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_277; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_278; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_279; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_280; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_281; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_282; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_283; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_284; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_285; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_286; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_287; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_288; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_289; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_290; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_291; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_292; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_293; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_294; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_295; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_296; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_297; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_298; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_299; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_300; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_301; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_302; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_303; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_304; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_305; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_306; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_307; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_308; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_309; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_310; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_311; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_312; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_313; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_314; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_315; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_316; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_317; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_318; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_319; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_320; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_321; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_322; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_323; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_324; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_325; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_326; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_327; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_328; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_329; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_330; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_331; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_332; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_333; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_334; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_335; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_336; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_337; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_338; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_339; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_340; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_341; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_342; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_343; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_344; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_345; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_346; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_347; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_348; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_349; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_350; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_351; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_352; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_353; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_354; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_355; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_356; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_357; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_358; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_359; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_360; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_361; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_362; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_363; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_364; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_365; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_366; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_367; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_368; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_369; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_370; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_371; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_372; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_373; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_374; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_375; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_376; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_377; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_378; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_379; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_380; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_381; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_382; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_383; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_384; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_385; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_386; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_387; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_388; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_389; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_390; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_391; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_392; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_393; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_394; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_395; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_396; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_397; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_398; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_399; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_400; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_401; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_402; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_403; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_404; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_405; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_406; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_407; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_408; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_409; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_410; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_411; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_412; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_413; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_414; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_415; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_416; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_417; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_418; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_419; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_420; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_421; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_422; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_423; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_424; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_425; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_426; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_427; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_428; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_429; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_430; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_431; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_432; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_433; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_434; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_435; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_436; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_437; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_438; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_439; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_440; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_441; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_442; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_443; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_444; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_445; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_446; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_447; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_448; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_449; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_450; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_451; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_452; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_453; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_454; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_455; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_456; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_457; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_458; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_459; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_460; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_461; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_462; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_463; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_464; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_465; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_466; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_467; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_468; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_469; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_470; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_471; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_472; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_473; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_474; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_475; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_476; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_477; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_478; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_479; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_480; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_481; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_482; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_483; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_484; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_485; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_486; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_487; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_488; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_489; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_490; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_491; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_492; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_493; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_494; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_495; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_496; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_497; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_498; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_499; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_500; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_501; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_502; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_503; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_504; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_505; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_506; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_507; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_508; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_509; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_510; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_511; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_512; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_513; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_514; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_515; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_516; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_517; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_518; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_519; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_520; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_521; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_522; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_523; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_524; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_525; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_526; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_527; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_528; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_529; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_530; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_531; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_532; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_533; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_534; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_535; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_536; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_537; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_538; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_539; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_540; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_541; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_542; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_543; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_544; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_545; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_546; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_547; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_548; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_549; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_550; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_551; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_552; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_553; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_554; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_555; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_556; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_557; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_558; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_559; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_560; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_561; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_562; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_563; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_564; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_565; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_566; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_567; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_568; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_569; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_570; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_571; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_572; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_573; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_574; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_575; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_576; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_577; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_578; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_579; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_580; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_581; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_582; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_583; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_584; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_585; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_586; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_587; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_588; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_589; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_590; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_591; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_592; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_593; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_594; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_595; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_596; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_597; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_598; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_599; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_600; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_601; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_602; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_603; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_604; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_605; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_606; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_607; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_608; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_609; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_610; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_611; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_612; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_613; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_614; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_615; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_616; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_617; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_618; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_619; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_620; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_621; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_622; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_623; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_624; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_625; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_626; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_627; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_628; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_629; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_630; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_631; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_632; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_633; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_634; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_635; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_636; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_637; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_638; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_639; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_640; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_641; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_642; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_643; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_644; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_645; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_646; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_647; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_648; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_649; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_650; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_651; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_652; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_653; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_654; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_655; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_656; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_657; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_658; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_659; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_660; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_661; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_662; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_663; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_664; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_665; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_666; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_667; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_668; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_669; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_670; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_671; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_672; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_673; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_674; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_675; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_676; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_677; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_678; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_679; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_680; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_681; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_682; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_683; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_684; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_685; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_686; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_687; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_688; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_689; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_690; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_691; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_692; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_693; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_694; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_695; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_696; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_697; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_698; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_699; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_700; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_701; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_702; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_703; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_704; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_705; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_706; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_707; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_708; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_709; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_710; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_711; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_712; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_713; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_714; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_715; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_716; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_717; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_718; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_719; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_720; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_721; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_722; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_723; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_724; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_725; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_726; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_727; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_728; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_729; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_730; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_731; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_732; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_733; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_734; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_735; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_736; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_737; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_738; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_739; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_740; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_741; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_742; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_743; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_744; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_745; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_746; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_747; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_748; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_749; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_750; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_751; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_752; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_753; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_754; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_755; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_756; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_757; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_758; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_759; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_760; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_761; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_762; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_763; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_764; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_765; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_766; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_767; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_768; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_769; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_770; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_771; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_772; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_773; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_774; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_775; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_776; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_777; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_778; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_779; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_780; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_781; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_782; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_783; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_784; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_785; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_786; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_787; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_788; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_789; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_790; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_791; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_792; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_793; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_794; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_795; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_796; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_797; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_798; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_799; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_800; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_801; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_802; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_803; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_804; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_805; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_806; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_807; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_808; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_809; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_810; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_811; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_812; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_813; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_814; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_815; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_816; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_817; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_818; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_819; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_820; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_821; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_822; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_823; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_824; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_825; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_826; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_827; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_828; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_829; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_830; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_831; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_832; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_833; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_834; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_835; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_836; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_837; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_838; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_839; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_840; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_841; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_842; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_843; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_844; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_845; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_846; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_847; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_848; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_849; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_850; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_851; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_852; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_853; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_854; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_855; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_856; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_857; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_858; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_859; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_860; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_861; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_862; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_863; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_864; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_865; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_866; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_867; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_868; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_869; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_870; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_871; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_872; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_873; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_874; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_875; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_876; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_877; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_878; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_879; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_880; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_881; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_882; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_883; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_884; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_885; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_886; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_887; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_888; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_889; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_890; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_891; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_892; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_893; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_894; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_895; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_896; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_897; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_898; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_899; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_900; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_901; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_902; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_903; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_904; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_905; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_906; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_907; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_908; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_909; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_910; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_911; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_912; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_913; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_914; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_915; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_916; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_917; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_918; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_919; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_920; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_921; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_922; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_923; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_924; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_925; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_926; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_927; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_928; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_929; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_930; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_931; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_932; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_933; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_934; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_935; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_936; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_937; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_938; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_939; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_940; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_941; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_942; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_943; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_944; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_945; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_946; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_947; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_948; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_949; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_950; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_951; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_952; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_953; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_954; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_955; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_956; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_957; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_958; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_959; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_960; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_961; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_962; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_963; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_964; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_965; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_966; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_967; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_968; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_969; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_970; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_971; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_972; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_973; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_974; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_975; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_976; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_977; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_978; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_979; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_980; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_981; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_982; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_983; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_984; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_985; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_986; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_987; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_988; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_989; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_990; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_991; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_992; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_993; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_994; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_995; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_996; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_997; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_998; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_999; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1000; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1001; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1002; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1003; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1004; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1005; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1006; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1007; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1008; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1009; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1010; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1011; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1012; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1013; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1014; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1015; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1016; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1017; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1018; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1019; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1020; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1021; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1022; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1023; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1024; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1025; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1026; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1027; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1028; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1029; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1030; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1031; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1032; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1033; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1034; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1035; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1036; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1037; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1038; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1039; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1040; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1041; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1042; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1043; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1044; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1045; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1046; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1047; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1048; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1049; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1050; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1051; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1052; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1053; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1054; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1055; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1056; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1057; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1058; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1059; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1060; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1061; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1062; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1063; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1064; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1065; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1066; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1067; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1068; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1069; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1070; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1071; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1072; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1073; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1074; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1075; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1076; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1077; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1078; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1079; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1080; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1081; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1082; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1083; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1084; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1085; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1086; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1087; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1088; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1089; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1090; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1091; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1092; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1093; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1094; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1095; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1096; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1097; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1098; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1099; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1100; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1101; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1102; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1103; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1104; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1105; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1106; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1107; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1108; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1109; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1110; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1111; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1112; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1113; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1114; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1115; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1116; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1117; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1118; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1119; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1120; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1121; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1122; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1123; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1124; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1125; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1126; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1127; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1128; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1129; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1130; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1131; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1132; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1133; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1134; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1135; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1136; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1137; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1138; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1139; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1140; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1141; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1142; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1143; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1144; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1145; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1146; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1147; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1148; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1149; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1150; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1151; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1152; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1153; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1154; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1155; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1156; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1157; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1158; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1159; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1160; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1161; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1162; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1163; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1164; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1165; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1166; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1167; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1168; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1169; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1170; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1171; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1172; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1173; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1174; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1175; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1176; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1177; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1178; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1179; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1180; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1181; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1182; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1183; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1184; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1185; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1186; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1187; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1188; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1189; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1190; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1191; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1192; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1193; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1194; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1195; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1196; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1197; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1198; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1199; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1200; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1201; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1202; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1203; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1204; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1205; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1206; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1207; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1208; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1209; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1210; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1211; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1212; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1213; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1214; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1215; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1216; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1217; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1218; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1219; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1220; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1221; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1222; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1223; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1224; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1225; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1226; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1227; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1228; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1229; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1230; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1231; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1232; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1233; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1234; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1235; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1236; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1237; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1238; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1239; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1240; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1241; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1242; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1243; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1244; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1245; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1246; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1247; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1248; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1249; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1250; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1251; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1252; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1253; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1254; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1255; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1256; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1257; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1258; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1259; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1260; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1261; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1262; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1263; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1264; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1265; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1266; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1267; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1268; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1269; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1270; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1271; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1272; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1273; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1274; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1275; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1276; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1277; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1278; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1279; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1280; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1281; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1282; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1283; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1284; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1285; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1286; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1287; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1288; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1289; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1290; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1291; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1292; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1293; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1294; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1295; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1296; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1297; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1298; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1299; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1300; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1301; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1302; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1303; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1304; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1305; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1306; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1307; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1308; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1309; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1310; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1311; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1312; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1313; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1314; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1315; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1316; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1317; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1318; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1319; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1320; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1321; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1322; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1323; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1324; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1325; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1326; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1327; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1328; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1329; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1330; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1331; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1332; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1333; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1334; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1335; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1336; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1337; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1338; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1339; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1340; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1341; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1342; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1343; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1344; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1345; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1346; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1347; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1348; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1349; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1350; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1351; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1352; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1353; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1354; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1355; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1356; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1357; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1358; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1359; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1360; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1361; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1362; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1363; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1364; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1365; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1366; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1367; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1368; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1369; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1370; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1371; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1372; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1373; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1374; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1375; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1376; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1377; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1378; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1379; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1380; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1381; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1382; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1383; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1384; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1385; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1386; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1387; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1388; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1389; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1390; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1391; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1392; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1393; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1394; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1395; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1396; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1397; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1398; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1399; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1400; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1401; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1402; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1403; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1404; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1405; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1406; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1407; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1408; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1409; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1410; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1411; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1412; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1413; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1414; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1415; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1416; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1417; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1418; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1419; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1420; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1421; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1422; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1423; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1424; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1425; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1426; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1427; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1428; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1429; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1430; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1431; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1432; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1433; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1434; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1435; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1436; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1437; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1438; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1439; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1440; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1441; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1442; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1443; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1444; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1445; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1446; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1447; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1448; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1449; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1450; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1451; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1452; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1453; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1454; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1455; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1456; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1457; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1458; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1459; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1460; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1461; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1462; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1463; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1464; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1465; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1466; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1467; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1468; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1469; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1470; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1471; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1472; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1473; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1474; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1475; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1476; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1477; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1478; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1479; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1480; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1481; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1482; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1483; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1484; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1485; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1486; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1487; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1488; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1489; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1490; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1491; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1492; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1493; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1494; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1495; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1496; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1497; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1498; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1499; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1500; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1501; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1502; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1503; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1504; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1505; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1506; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1507; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1508; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1509; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1510; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1511; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1512; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1513; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1514; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1515; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1516; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1517; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1518; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1519; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1520; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1521; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1522; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1523; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1524; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1525; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1526; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1527; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1528; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1529; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1530; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1531; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1532; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1533; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1534; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1535; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1536; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1537; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1538; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1539; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1540; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1541; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1542; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1543; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1544; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1545; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1546; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1547; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1548; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1549; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1550; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1551; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1552; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1553; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1554; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1555; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1556; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1557; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1558; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1559; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1560; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1561; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1562; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1563; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1564; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1565; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1566; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1567; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1568; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1569; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1570; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1571; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1572; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1573; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1574; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1575; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1576; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1577; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1578; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1579; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1580; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1581; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1582; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1583; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1584; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1585; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1586; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1587; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1588; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1589; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1590; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1591; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1592; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1593; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1594; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1595; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1596; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1597; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1598; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1599; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1600; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1601; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1602; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1603; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1604; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1605; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1606; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1607; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1608; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1609; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1610; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1611; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1612; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1613; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1614; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1615; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1616; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1617; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1618; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1619; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1620; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1621; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1622; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1623; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1624; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1625; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1626; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1627; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1628; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1629; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1630; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1631; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1632; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1633; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1634; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1635; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1636; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1637; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1638; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1639; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1640; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1641; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1642; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1643; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1644; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1645; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1646; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1647; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1648; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1649; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1650; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1651; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1652; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1653; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1654; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1655; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1656; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1657; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1658; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1659; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1660; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1661; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1662; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1663; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1664; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1665; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1666; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1667; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1668; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1669; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1670; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1671; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1672; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1673; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1674; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1675; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1676; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1677; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1678; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1679; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1680; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1681; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1682; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1683; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1684; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1685; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1686; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1687; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1688; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1689; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1690; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1691; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1692; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1693; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1694; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1695; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1696; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1697; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1698; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1699; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1700; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1701; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1702; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1703; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1704; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1705; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1706; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1707; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1708; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1709; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1710; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1711; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1712; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1713; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1714; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1715; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1716; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1717; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1718; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1719; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1720; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1721; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1722; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1723; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1724; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1725; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1726; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1727; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1728; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1729; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1730; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1731; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1732; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1733; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1734; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1735; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1736; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1737; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1738; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1739; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1740; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1741; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1742; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1743; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1744; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1745; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1746; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1747; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1748; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1749; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1750; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1751; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1752; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1753; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1754; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1755; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1756; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1757; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1758; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1759; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1760; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1761; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1762; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1763; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1764; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1765; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1766; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1767; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1768; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1769; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1770; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1771; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1772; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1773; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1774; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1775; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1776; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1777; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1778; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1779; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1780; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1781; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1782; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1783; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1784; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1785; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1786; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1787; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1788; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1789; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1790; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1791; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1792; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1793; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1794; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1795; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1796; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1797; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1798; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1799; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1800; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1801; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1802; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1803; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1804; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1805; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1806; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1807; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1808; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1809; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1810; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1811; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1812; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1813; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1814; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1815; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1816; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1817; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1818; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1819; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1820; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1821; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1822; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1823; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1824; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1825; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1826; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1827; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1828; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1829; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1830; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1831; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1832; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1833; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1834; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1835; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1836; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1837; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1838; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1839; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1840; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1841; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1842; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1843; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1844; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1845; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1846; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1847; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1848; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1849; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1850; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1851; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1852; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1853; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1854; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1855; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1856; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1857; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1858; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1859; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1860; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1861; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1862; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1863; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1864; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1865; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1866; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1867; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1868; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1869; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1870; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1871; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1872; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1873; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1874; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1875; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1876; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1877; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1878; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1879; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1880; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1881; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1882; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1883; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1884; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1885; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1886; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1887; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1888; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1889; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1890; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1891; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1892; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1893; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1894; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1895; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1896; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1897; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1898; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1899; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1900; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1901; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1902; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1903; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1904; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1905; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1906; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1907; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1908; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1909; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1910; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1911; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1912; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1913; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1914; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1915; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1916; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1917; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1918; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1919; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1920; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1921; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1922; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1923; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1924; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1925; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1926; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1927; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1928; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1929; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1930; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1931; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1932; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1933; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1934; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1935; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1936; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1937; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1938; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1939; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1940; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1941; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1942; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1943; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1944; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1945; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1946; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1947; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1948; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1949; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1950; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1951; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1952; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1953; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1954; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1955; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1956; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1957; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1958; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1959; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1960; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1961; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1962; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1963; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1964; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1965; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1966; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1967; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1968; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1969; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1970; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1971; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1972; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1973; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1974; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1975; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1976; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1977; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1978; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1979; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1980; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1981; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1982; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1983; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1984; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1985; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1986; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1987; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1988; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1989; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1990; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1991; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1992; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1993; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1994; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1995; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1996; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1997; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1998; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_1999; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2000; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2001; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2002; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2003; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2004; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2005; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2006; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2007; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2008; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2009; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2010; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2011; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2012; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2013; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2014; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2015; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2016; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2017; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2018; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2019; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2020; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2021; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2022; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2023; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2024; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2025; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2026; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2027; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2028; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2029; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2030; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2031; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2032; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2033; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2034; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2035; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2036; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2037; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2038; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2039; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2040; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2041; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2042; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2043; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2044; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2045; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2046; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2047; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2048; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2049; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2050; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2051; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2052; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2053; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2054; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2055; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2056; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2057; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2058; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2059; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2060; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2061; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2062; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2063; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2064; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2065; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2066; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2067; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2068; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2069; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2070; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2071; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2072; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2073; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2074; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2075; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2076; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2077; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2078; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2079; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2080; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2081; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2082; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2083; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2084; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2085; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2086; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2087; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2088; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2089; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2090; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2091; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2092; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2093; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2094; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2095; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2096; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2097; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2098; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2099; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2100; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2101; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2102; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2103; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2104; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2105; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2106; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2107; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2108; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2109; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2110; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2111; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2112; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2113; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2114; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2115; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2116; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2117; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2118; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2119; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2120; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2121; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2122; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2123; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2124; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2125; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2126; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2127; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2128; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2129; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2130; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2131; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2132; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2133; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2134; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2135; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2136; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2137; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2138; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2139; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2140; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2141; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2142; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2143; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2144; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2145; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2146; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2147; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2148; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2149; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2150; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2151; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2152; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2153; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2154; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2155; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2156; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2157; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2158; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2159; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2160; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2161; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2162; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2163; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2164; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2165; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2166; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2167; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2168; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2169; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2170; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2171; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2172; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2173; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2174; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2175; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2176; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2177; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2178; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2179; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2180; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2181; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2182; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2183; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2184; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2185; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2186; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2187; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2188; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2189; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2190; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2191; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2192; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2193; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2194; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2195; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2196; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2197; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2198; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2199; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2200; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2201; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2202; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2203; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2204; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2205; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2206; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2207; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2208; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2209; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2210; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2211; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2212; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2213; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2214; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2215; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2216; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2217; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2218; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2219; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2220; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2221; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2222; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2223; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2224; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2225; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2226; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2227; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2228; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2229; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2230; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2231; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2232; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2233; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2234; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2235; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2236; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2237; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2238; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2239; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2240; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2241; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2242; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2243; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2244; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2245; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2246; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2247; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2248; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2249; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2250; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2251; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2252; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2253; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2254; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2255; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2256; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2257; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2258; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2259; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2260; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2261; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2262; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2263; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2264; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2265; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2266; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2267; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2268; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2269; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2270; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2271; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2272; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2273; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2274; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2275; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2276; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2277; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2278; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2279; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2280; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2281; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2282; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2283; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2284; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2285; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2286; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2287; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2288; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2289; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2290; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2291; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2292; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2293; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2294; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2295; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2296; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2297; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2298; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2299; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2300; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2301; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2302; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2303; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2304; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2305; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2306; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2307; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2308; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2309; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2310; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2311; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2312; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2313; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2314; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2315; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2316; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2317; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2318; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2319; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2320; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2321; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2322; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2323; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2324; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2325; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2326; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2327; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2328; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2329; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2330; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2331; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2332; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2333; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2334; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2335; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2336; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2337; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2338; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2339; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2340; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2341; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2342; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2343; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2344; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2345; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2346; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2347; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2348; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2349; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2350; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2351; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2352; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2353; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2354; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2355; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2356; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2357; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2358; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2359; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2360; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2361; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2362; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2363; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2364; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2365; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2366; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2367; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2368; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2369; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2370; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2371; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2372; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2373; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2374; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2375; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2376; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2377; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2378; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2379; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2380; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2381; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2382; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2383; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2384; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2385; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2386; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2387; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2388; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2389; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2390; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2391; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2392; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2393; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2394; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2395; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2396; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2397; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2398; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2399; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2400; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2401; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2402; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2403; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2404; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2405; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2406; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2407; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2408; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2409; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2410; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2411; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2412; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2413; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2414; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2415; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2416; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2417; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2418; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2419; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2420; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2421; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2422; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2423; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2424; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2425; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2426; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2427; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2428; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2429; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2430; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2431; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2432; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2433; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2434; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2435; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2436; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2437; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2438; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2439; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2440; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2441; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2442; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2443; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2444; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2445; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2446; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2447; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2448; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2449; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2450; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2451; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2452; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2453; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2454; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2455; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2456; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2457; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2458; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2459; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2460; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2461; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2462; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2463; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2464; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2465; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2466; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2467; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2468; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2469; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2470; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2471; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2472; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2473; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2474; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2475; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2476; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2477; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2478; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2479; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2480; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2481; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2482; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2483; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2484; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2485; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2486; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2487; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2488; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2489; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2490; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2491; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2492; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2493; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2494; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2495; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2496; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2497; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2498; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2499; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2500; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2501; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2502; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2503; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2504; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2505; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2506; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2507; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2508; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2509; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2510; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2511; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2512; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2513; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2514; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2515; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2516; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2517; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2518; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2519; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2520; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2521; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2522; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2523; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2524; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2525; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2526; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2527; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2528; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2529; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2530; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2531; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2532; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2533; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2534; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2535; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2536; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2537; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2538; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2539; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2540; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2541; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2542; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2543; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2544; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2545; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2546; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2547; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2548; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2549; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2550; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2551; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2552; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2553; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2554; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2555; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2556; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2557; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2558; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2559; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2560; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2561; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2562; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2563; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2564; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2565; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2566; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2567; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2568; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2569; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2570; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2571; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2572; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2573; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2574; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2575; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2576; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2577; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2578; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2579; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2580; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2581; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2582; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2583; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2584; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2585; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2586; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2587; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2588; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2589; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2590; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2591; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2592; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2593; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2594; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2595; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2596; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2597; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2598; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2599; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2600; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2601; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2602; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2603; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2604; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2605; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2606; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2607; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2608; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2609; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2610; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2611; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2612; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2613; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2614; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2615; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2616; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2617; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2618; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2619; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2620; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2621; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2622; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2623; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2624; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2625; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2626; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2627; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2628; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2629; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2630; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2631; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2632; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2633; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2634; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2635; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2636; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2637; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2638; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2639; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2640; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2641; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2642; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2643; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2644; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2645; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2646; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2647; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2648; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2649; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2650; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2651; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2652; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2653; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2654; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2655; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2656; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2657; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2658; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2659; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2660; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2661; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2662; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2663; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2664; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2665; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2666; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2667; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2668; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2669; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2670; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2671; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2672; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2673; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2674; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2675; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2676; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2677; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2678; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2679; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2680; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2681; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2682; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2683; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2684; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2685; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2686; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2687; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2688; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2689; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2690; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2691; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2692; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2693; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2694; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2695; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2696; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2697; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2698; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2699; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2700; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2701; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2702; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2703; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2704; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2705; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2706; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2707; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2708; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2709; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2710; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2711; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2712; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2713; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2714; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2715; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2716; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2717; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2718; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2719; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2720; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2721; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2722; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2723; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2724; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2725; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2726; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2727; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2728; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2729; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2730; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2731; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2732; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2733; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2734; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2735; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2736; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2737; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2738; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2739; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2740; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2741; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2742; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2743; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2744; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2745; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2746; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2747; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2748; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2749; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2750; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2751; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2752; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2753; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2754; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2755; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2756; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2757; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2758; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2759; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2760; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2761; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2762; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2763; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2764; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2765; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2766; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2767; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2768; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2769; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2770; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2771; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2772; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2773; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2774; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2775; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2776; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2777; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2778; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2779; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2780; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2781; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2782; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2783; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2784; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2785; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2786; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2787; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2788; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2789; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2790; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2791; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2792; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2793; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2794; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2795; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2796; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2797; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2798; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2799; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2800; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2801; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2802; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2803; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2804; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2805; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2806; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2807; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2808; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2809; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2810; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2811; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2812; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2813; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2814; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2815; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2816; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2817; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2818; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2819; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2820; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2821; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2822; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2823; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2824; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2825; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2826; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2827; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2828; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2829; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2830; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2831; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2832; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2833; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2834; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2835; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2836; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2837; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2838; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2839; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2840; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2841; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2842; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2843; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2844; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2845; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2846; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2847; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2848; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2849; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2850; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2851; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2852; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2853; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2854; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2855; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2856; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2857; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2858; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2859; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2860; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2861; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2862; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2863; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2864; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2865; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2866; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2867; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2868; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2869; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2870; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2871; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2872; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2873; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2874; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2875; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2876; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2877; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2878; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2879; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2880; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2881; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2882; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2883; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2884; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2885; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2886; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2887; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2888; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2889; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2890; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2891; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2892; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2893; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2894; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2895; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2896; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2897; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2898; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2899; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2900; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2901; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2902; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2903; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2904; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2905; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2906; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2907; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2908; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2909; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2910; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2911; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2912; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2913; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2914; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2915; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2916; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2917; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2918; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2919; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2920; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2921; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2922; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2923; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2924; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2925; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2926; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2927; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2928; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2929; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2930; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2931; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2932; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2933; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2934; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2935; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2936; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2937; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2938; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2939; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2940; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2941; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2942; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2943; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2944; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2945; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2946; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2947; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2948; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2949; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2950; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2951; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2952; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2953; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2954; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2955; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2956; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2957; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2958; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2959; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2960; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2961; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2962; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2963; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2964; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2965; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2966; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2967; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2968; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2969; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2970; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2971; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2972; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2973; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2974; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2975; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2976; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2977; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2978; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2979; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2980; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2981; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2982; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2983; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2984; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2985; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2986; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2987; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2988; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2989; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2990; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2991; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2992; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2993; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2994; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2995; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2996; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2997; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2998; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_2999; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3000; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3001; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3002; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3003; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3004; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3005; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3006; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3007; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3008; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3009; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3010; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3011; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3012; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3013; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3014; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3015; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3016; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3017; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3018; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3019; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3020; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3021; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3022; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3023; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3024; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3025; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3026; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3027; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3028; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3029; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3030; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3031; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3032; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3033; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3034; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3035; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3036; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3037; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3038; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3039; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3040; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3041; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3042; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3043; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3044; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3045; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3046; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3047; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3048; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3049; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3050; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3051; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3052; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3053; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3054; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3055; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3056; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3057; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3058; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3059; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3060; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3061; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3062; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3063; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3064; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3065; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3066; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3067; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3068; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3069; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3070; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3071; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3072; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3073; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3074; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3075; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3076; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3077; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3078; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3079; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3080; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3081; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3082; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3083; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3084; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3085; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3086; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3087; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3088; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3089; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3090; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3091; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3092; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3093; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3094; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3095; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3096; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3097; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3098; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3099; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3100; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3101; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3102; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3103; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3104; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3105; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3106; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3107; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3108; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3109; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3110; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3111; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3112; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3113; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3114; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3115; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3116; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3117; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3118; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3119; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3120; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3121; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3122; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3123; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3124; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3125; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3126; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3127; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3128; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3129; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3130; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3131; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3132; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3133; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3134; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3135; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3136; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3137; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3138; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3139; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3140; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3141; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3142; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3143; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3144; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3145; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3146; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3147; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3148; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3149; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3150; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3151; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3152; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3153; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3154; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3155; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3156; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3157; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3158; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3159; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3160; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3161; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3162; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3163; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3164; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3165; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3166; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3167; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3168; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3169; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3170; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3171; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3172; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3173; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3174; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3175; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3176; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3177; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3178; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3179; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3180; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3181; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3182; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3183; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3184; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3185; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3186; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3187; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3188; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3189; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3190; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3191; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3192; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3193; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3194; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3195; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3196; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3197; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3198; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3199; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3200; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3201; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3202; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3203; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3204; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3205; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3206; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3207; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3208; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3209; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3210; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3211; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3212; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3213; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3214; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3215; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3216; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3217; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3218; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3219; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3220; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3221; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3222; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3223; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3224; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3225; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3226; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3227; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3228; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3229; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3230; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3231; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3232; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3233; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3234; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3235; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3236; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3237; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3238; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3239; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3240; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3241; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3242; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3243; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3244; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3245; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3246; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3247; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3248; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3249; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3250; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3251; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3252; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3253; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3254; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3255; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3256; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3257; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3258; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3259; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3260; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3261; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3262; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3263; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3264; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3265; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3266; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3267; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3268; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3269; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3270; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3271; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3272; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3273; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3274; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3275; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3276; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3277; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3278; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3279; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3280; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3281; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3282; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3283; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3284; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3285; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3286; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3287; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3288; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3289; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3290; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3291; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3292; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3293; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3294; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3295; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3296; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3297; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3298; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3299; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3300; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3301; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3302; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3303; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3304; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3305; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3306; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3307; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3308; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3309; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3310; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3311; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3312; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3313; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3314; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3315; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3316; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3317; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3318; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3319; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3320; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3321; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3322; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3323; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3324; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3325; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3326; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3327; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3328; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3329; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3330; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3331; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3332; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3333; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3334; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3335; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3336; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3337; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3338; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3339; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3340; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3341; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3342; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3343; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3344; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3345; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3346; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3347; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3348; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3349; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3350; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3351; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3352; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3353; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3354; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3355; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3356; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3357; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3358; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3359; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3360; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3361; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3362; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3363; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3364; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3365; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3366; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3367; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3368; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3369; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3370; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3371; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3372; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3373; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3374; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3375; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3376; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3377; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3378; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3379; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3380; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3381; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3382; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3383; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3384; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3385; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3386; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3387; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3388; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3389; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3390; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3391; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3392; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3393; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3394; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3395; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3396; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3397; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3398; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3399; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3400; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3401; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3402; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3403; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3404; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3405; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3406; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3407; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3408; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3409; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3410; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3411; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3412; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3413; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3414; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3415; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3416; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3417; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3418; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3419; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3420; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3421; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3422; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3423; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3424; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3425; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3426; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3427; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3428; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3429; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3430; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3431; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3432; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3433; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3434; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3435; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3436; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3437; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3438; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3439; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3440; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3441; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3442; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3443; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3444; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3445; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3446; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3447; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3448; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3449; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3450; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3451; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3452; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3453; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3454; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3455; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3456; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3457; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3458; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3459; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3460; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3461; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3462; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3463; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3464; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3465; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3466; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3467; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3468; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3469; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3470; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3471; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3472; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3473; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3474; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3475; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3476; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3477; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3478; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3479; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3480; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3481; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3482; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3483; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3484; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3485; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3486; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3487; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3488; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3489; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3490; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3491; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3492; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3493; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3494; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3495; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3496; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3497; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3498; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3499; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3500; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3501; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3502; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3503; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3504; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3505; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3506; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3507; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3508; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3509; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3510; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3511; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3512; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3513; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3514; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3515; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3516; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3517; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3518; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3519; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3520; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3521; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3522; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3523; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3524; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3525; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3526; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3527; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3528; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3529; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3530; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3531; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3532; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3533; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3534; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3535; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3536; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3537; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3538; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3539; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3540; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3541; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3542; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3543; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3544; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3545; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3546; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3547; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3548; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3549; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3550; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3551; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3552; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3553; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3554; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3555; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3556; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3557; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3558; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3559; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3560; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3561; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3562; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3563; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3564; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3565; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3566; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3567; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3568; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3569; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3570; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3571; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3572; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3573; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3574; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3575; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3576; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3577; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3578; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3579; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3580; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3581; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3582; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3583; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3584; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3585; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3586; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3587; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3588; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3589; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3590; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3591; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3592; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3593; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3594; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3595; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3596; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3597; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3598; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3599; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3600; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3601; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3602; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3603; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3604; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3605; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3606; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3607; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3608; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3609; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3610; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3611; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3612; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3613; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3614; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3615; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3616; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3617; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3618; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3619; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3620; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3621; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3622; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3623; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3624; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3625; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3626; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3627; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3628; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3629; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3630; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3631; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3632; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3633; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3634; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3635; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3636; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3637; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3638; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3639; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3640; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3641; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3642; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3643; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3644; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3645; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3646; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3647; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3648; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3649; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3650; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3651; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3652; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3653; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3654; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3655; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3656; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3657; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3658; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3659; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3660; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3661; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3662; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3663; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3664; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3665; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3666; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3667; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3668; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3669; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3670; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3671; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3672; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3673; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3674; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3675; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3676; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3677; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3678; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3679; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3680; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3681; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3682; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3683; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3684; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3685; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3686; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3687; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3688; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3689; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3690; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3691; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3692; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3693; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3694; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3695; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3696; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3697; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3698; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3699; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3700; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3701; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3702; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3703; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3704; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3705; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3706; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3707; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3708; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3709; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3710; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3711; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3712; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3713; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3714; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3715; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3716; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3717; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3718; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3719; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3720; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3721; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3722; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3723; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3724; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3725; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3726; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3727; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3728; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3729; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3730; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3731; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3732; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3733; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3734; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3735; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3736; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3737; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3738; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3739; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3740; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3741; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3742; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3743; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3744; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3745; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3746; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3747; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3748; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3749; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3750; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3751; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3752; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3753; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3754; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3755; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3756; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3757; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3758; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3759; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3760; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3761; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3762; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3763; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3764; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3765; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3766; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3767; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3768; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3769; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3770; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3771; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3772; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3773; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3774; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3775; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3776; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3777; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3778; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3779; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3780; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3781; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3782; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3783; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3784; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3785; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3786; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3787; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3788; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3789; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3790; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3791; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3792; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3793; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3794; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3795; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3796; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3797; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3798; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3799; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3800; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3801; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3802; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3803; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3804; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3805; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3806; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3807; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3808; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3809; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3810; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3811; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3812; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3813; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3814; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3815; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3816; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3817; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3818; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3819; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3820; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3821; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3822; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3823; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3824; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3825; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3826; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3827; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3828; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3829; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3830; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3831; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3832; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3833; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3834; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3835; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3836; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3837; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3838; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3839; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3840; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3841; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3842; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3843; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3844; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3845; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3846; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3847; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3848; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3849; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3850; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3851; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3852; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3853; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3854; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3855; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3856; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3857; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3858; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3859; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3860; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3861; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3862; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3863; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3864; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3865; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3866; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3867; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3868; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3869; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3870; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3871; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3872; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3873; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3874; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3875; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3876; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3877; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3878; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3879; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3880; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3881; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3882; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3883; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3884; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3885; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3886; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3887; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3888; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3889; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3890; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3891; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3892; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3893; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3894; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3895; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3896; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3897; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3898; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3899; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3900; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3901; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3902; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3903; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3904; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3905; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3906; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3907; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3908; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3909; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3910; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3911; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3912; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3913; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3914; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3915; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3916; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3917; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3918; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3919; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3920; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3921; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3922; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3923; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3924; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3925; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3926; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3927; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3928; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3929; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3930; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3931; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3932; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3933; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3934; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3935; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3936; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3937; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3938; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3939; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3940; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3941; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3942; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3943; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3944; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3945; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3946; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3947; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3948; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3949; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3950; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3951; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3952; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3953; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3954; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3955; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3956; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3957; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3958; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3959; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3960; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3961; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3962; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3963; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3964; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3965; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3966; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3967; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3968; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3969; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3970; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3971; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3972; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3973; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3974; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3975; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3976; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3977; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3978; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3979; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3980; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3981; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3982; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3983; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3984; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3985; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3986; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3987; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3988; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3989; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3990; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3991; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3992; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3993; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3994; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3995; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3996; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3997; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3998; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_3999; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4000; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4001; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4002; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4003; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4004; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4005; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4006; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4007; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4008; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4009; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4010; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4011; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4012; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4013; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4014; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4015; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4016; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4017; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4018; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4019; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4020; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4021; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4022; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4023; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4024; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4025; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4026; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4027; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4028; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4029; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4030; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4031; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4032; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4033; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4034; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4035; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4036; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4037; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4038; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4039; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4040; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4041; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4042; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4043; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4044; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4045; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4046; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4047; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4048; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4049; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4050; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4051; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4052; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4053; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4054; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4055; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4056; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4057; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4058; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4059; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4060; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4061; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4062; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4063; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4064; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4065; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4066; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4067; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4068; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4069; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4070; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4071; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4072; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4073; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4074; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4075; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4076; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4077; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4078; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4079; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4080; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4081; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4082; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4083; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4084; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4085; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4086; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4087; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4088; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4089; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4090; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4091; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4092; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4093; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4094; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4095; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4096; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4097; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4098; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4099; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4100; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4101; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4102; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4103; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4104; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4105; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4106; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4107; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4108; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4109; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4110; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4111; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4112; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4113; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4114; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4115; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4116; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4117; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4118; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4119; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4120; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4121; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4122; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4123; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4124; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4125; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4126; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4127; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4128; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4129; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4130; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4131; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4132; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4133; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4134; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4135; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4136; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4137; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4138; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4139; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4140; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4141; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4142; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4143; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4144; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4145; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4146; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4147; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4148; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4149; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4150; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4151; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4152; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4153; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4154; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4155; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4156; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4157; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4158; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4159; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4160; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4161; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4162; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4163; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4164; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4165; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4166; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4167; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4168; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4169; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4170; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4171; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4172; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4173; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4174; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4175; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4176; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4177; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4178; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4179; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4180; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4181; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4182; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4183; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4184; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4185; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4186; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4187; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4188; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4189; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4190; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4191; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4192; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4193; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4194; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4195; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4196; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4197; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4198; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4199; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4200; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4201; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4202; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4203; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4204; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4205; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4206; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4207; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4208; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4209; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4210; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4211; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4212; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4213; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4214; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4215; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4216; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4217; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4218; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4219; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4220; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4221; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4222; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4223; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4224; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4225; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4226; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4227; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4228; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4229; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4230; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4231; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4232; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4233; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4234; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4235; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4236; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4237; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4238; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4239; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4240; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4241; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4242; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4243; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4244; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4245; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4246; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4247; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4248; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4249; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4250; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4251; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4252; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4253; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4254; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4255; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4256; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4257; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4258; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4259; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4260; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4261; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4262; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4263; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4264; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4265; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4266; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4267; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4268; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4269; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4270; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4271; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4272; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4273; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4274; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4275; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4276; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4277; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4278; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4279; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4280; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4281; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4282; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4283; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4284; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4285; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4286; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4287; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4288; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4289; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4290; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4291; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4292; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4293; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4294; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4295; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4296; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4297; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4298; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4299; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4300; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4301; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4302; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4303; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4304; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4305; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4306; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4307; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4308; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4309; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4310; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4311; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4312; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4313; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4314; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4315; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4316; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4317; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4318; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4319; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4320; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4321; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4322; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4323; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4324; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4325; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4326; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4327; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4328; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4329; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4330; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4331; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4332; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4333; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4334; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4335; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4336; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4337; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4338; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4339; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4340; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4341; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4342; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4343; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4344; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4345; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4346; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4347; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4348; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4349; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4350; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4351; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4352; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4353; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4354; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4355; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4356; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4357; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4358; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4359; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4360; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4361; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4362; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4363; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4364; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4365; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4366; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4367; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4368; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4369; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4370; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4371; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4372; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4373; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4374; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4375; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4376; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4377; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4378; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4379; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4380; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4381; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4382; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4383; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4384; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4385; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4386; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4387; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4388; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4389; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4390; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4391; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4392; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4393; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4394; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4395; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4396; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4397; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4398; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4399; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4400; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4401; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4402; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4403; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4404; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4405; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4406; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4407; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4408; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4409; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4410; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4411; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4412; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4413; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4414; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4415; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4416; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4417; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4418; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4419; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4420; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4421; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4422; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4423; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4424; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4425; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4426; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4427; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4428; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4429; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4430; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4431; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4432; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4433; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4434; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4435; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4436; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4437; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4438; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4439; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4440; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4441; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4442; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4443; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4444; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4445; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4446; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4447; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4448; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4449; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4450; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4451; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4452; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4453; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4454; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4455; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4456; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4457; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4458; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4459; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4460; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4461; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4462; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4463; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4464; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4465; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4466; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4467; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4468; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4469; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4470; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4471; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4472; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4473; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4474; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4475; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4476; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4477; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4478; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4479; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4480; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4481; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4482; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4483; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4484; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4485; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4486; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4487; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4488; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4489; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4490; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4491; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4492; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4493; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4494; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4495; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4496; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4497; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4498; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4499; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4500; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4501; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4502; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4503; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4504; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4505; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4506; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4507; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4508; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4509; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4510; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4511; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4512; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4513; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4514; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4515; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4516; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4517; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4518; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4519; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4520; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4521; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4522; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4523; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4524; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4525; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4526; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4527; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4528; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4529; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4530; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4531; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4532; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4533; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4534; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4535; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4536; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4537; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4538; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4539; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4540; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4541; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4542; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4543; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4544; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4545; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4546; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4547; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4548; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4549; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4550; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4551; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4552; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4553; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4554; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4555; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4556; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4557; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4558; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4559; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4560; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4561; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4562; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4563; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4564; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4565; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4566; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4567; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4568; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4569; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4570; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4571; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4572; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4573; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4574; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4575; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4576; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4577; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4578; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4579; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4580; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4581; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4582; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4583; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4584; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4585; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4586; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4587; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4588; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4589; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4590; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4591; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4592; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4593; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4594; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4595; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4596; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4597; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4598; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4599; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4600; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4601; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4602; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4603; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4604; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4605; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4606; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4607; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4608; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4609; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4610; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4611; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4612; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4613; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4614; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4615; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4616; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4617; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4618; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4619; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4620; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4621; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4622; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4623; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4624; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4625; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4626; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4627; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4628; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4629; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4630; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4631; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4632; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4633; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4634; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4635; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4636; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4637; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4638; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4639; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4640; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4641; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4642; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4643; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4644; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4645; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4646; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4647; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4648; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4649; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4650; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4651; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4652; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4653; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4654; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4655; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4656; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4657; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4658; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4659; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4660; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4661; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4662; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4663; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4664; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4665; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4666; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4667; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4668; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4669; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4670; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4671; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4672; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4673; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4674; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4675; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4676; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4677; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4678; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4679; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4680; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4681; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4682; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4683; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4684; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4685; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4686; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4687; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4688; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4689; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4690; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4691; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4692; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4693; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4694; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4695; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4696; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4697; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4698; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4699; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4700; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4701; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4702; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4703; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4704; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4705; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4706; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4707; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4708; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4709; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4710; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4711; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4712; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4713; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4714; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4715; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4716; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4717; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4718; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4719; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4720; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4721; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4722; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4723; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4724; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4725; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4726; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4727; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4728; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4729; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4730; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4731; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4732; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4733; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4734; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4735; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4736; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4737; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4738; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4739; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4740; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4741; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4742; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4743; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4744; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4745; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4746; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4747; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4748; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4749; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4750; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4751; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4752; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4753; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4754; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4755; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4756; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4757; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4758; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4759; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4760; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4761; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4762; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4763; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4764; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4765; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4766; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4767; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4768; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4769; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4770; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4771; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4772; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4773; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4774; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4775; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4776; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4777; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4778; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4779; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4780; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4781; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4782; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4783; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4784; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4785; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4786; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4787; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4788; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4789; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4790; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4791; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4792; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4793; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4794; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4795; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4796; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4797; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4798; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4799; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4800; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4801; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4802; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4803; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4804; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4805; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4806; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4807; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4808; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4809; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4810; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4811; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4812; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4813; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4814; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4815; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4816; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4817; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4818; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4819; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4820; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4821; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4822; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4823; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4824; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4825; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4826; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4827; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4828; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4829; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4830; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4831; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4832; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4833; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4834; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4835; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4836; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4837; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4838; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4839; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4840; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4841; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4842; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4843; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4844; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4845; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4846; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4847; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4848; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4849; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4850; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4851; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4852; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4853; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4854; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4855; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4856; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4857; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4858; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4859; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4860; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4861; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4862; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4863; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4864; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4865; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4866; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4867; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4868; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4869; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4870; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4871; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4872; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4873; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4874; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4875; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4876; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4877; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4878; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4879; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4880; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4881; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4882; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4883; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4884; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4885; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4886; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4887; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4888; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4889; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4890; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4891; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4892; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4893; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4894; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4895; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4896; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4897; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4898; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4899; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4900; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4901; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4902; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4903; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4904; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4905; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4906; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4907; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4908; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4909; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4910; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4911; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4912; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4913; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4914; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4915; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4916; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4917; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4918; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4919; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4920; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4921; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4922; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4923; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4924; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4925; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4926; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4927; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4928; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4929; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4930; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4931; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4932; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4933; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4934; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4935; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4936; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4937; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4938; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4939; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4940; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4941; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4942; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4943; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4944; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4945; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4946; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4947; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4948; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4949; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4950; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4951; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4952; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4953; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4954; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4955; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4956; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4957; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4958; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4959; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4960; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4961; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4962; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4963; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4964; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4965; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4966; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4967; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4968; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4969; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4970; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4971; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4972; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4973; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4974; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4975; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4976; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4977; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4978; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4979; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4980; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4981; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4982; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4983; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4984; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4985; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4986; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4987; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4988; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4989; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4990; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4991; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4992; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4993; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4994; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4995; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4996; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4997; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4998; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_4999; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5000; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5001; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5002; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5003; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5004; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5005; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5006; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5007; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5008; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5009; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5010; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5011; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5012; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5013; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5014; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5015; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5016; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5017; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5018; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5019; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5020; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5021; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5022; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5023; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5024; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5025; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5026; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5027; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5028; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5029; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5030; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5031; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5032; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5033; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5034; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5035; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5036; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5037; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5038; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5039; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5040; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5041; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5042; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5043; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5044; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5045; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5046; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5047; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5048; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5049; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5050; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5051; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5052; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5053; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5054; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5055; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5056; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5057; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5058; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5059; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5060; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5061; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5062; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5063; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5064; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5065; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5066; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5067; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5068; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5069; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5070; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5071; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5072; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5073; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5074; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5075; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5076; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5077; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5078; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5079; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5080; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5081; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5082; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5083; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5084; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5085; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5086; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5087; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5088; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5089; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5090; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5091; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5092; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5093; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5094; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5095; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5096; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5097; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5098; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5099; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5100; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5101; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5102; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5103; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5104; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5105; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5106; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5107; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5108; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5109; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5110; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5111; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5112; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5113; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5114; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5115; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5116; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5117; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5118; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5119; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5120; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5121; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5122; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5123; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5124; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5125; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5126; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5127; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5128; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5129; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5130; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5131; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5132; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5133; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5134; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5135; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5136; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5137; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5138; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5139; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5140; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5141; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5142; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5143; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5144; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5145; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5146; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5147; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5148; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5149; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5150; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5151; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5152; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5153; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5154; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5155; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5156; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5157; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5158; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5159; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5160; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5161; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5162; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5163; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5164; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5165; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5166; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5167; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5168; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5169; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5170; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5171; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5172; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5173; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5174; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5175; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5176; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5177; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5178; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5179; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5180; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5181; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5182; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5183; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5184; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5185; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5186; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5187; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5188; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5189; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5190; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5191; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5192; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5193; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5194; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5195; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5196; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5197; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5198; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5199; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5200; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5201; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5202; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5203; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5204; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5205; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5206; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5207; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5208; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5209; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5210; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5211; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5212; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5213; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5214; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5215; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5216; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5217; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5218; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5219; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5220; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5221; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5222; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5223; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5224; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5225; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5226; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5227; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5228; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5229; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5230; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5231; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5232; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5233; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5234; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5235; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5236; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5237; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5238; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5239; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5240; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5241; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5242; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5243; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5244; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5245; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5246; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5247; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5248; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5249; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5250; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5251; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5252; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5253; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5254; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5255; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5256; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5257; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5258; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5259; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5260; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5261; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5262; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5263; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5264; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5265; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5266; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5267; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5268; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5269; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5270; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5271; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5272; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5273; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5274; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5275; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5276; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5277; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5278; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5279; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5280; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5281; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5282; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5283; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5284; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5285; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5286; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5287; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5288; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5289; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5290; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5291; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5292; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5293; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5294; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5295; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5296; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5297; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5298; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5299; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5300; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5301; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5302; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5303; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5304; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5305; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5306; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5307; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5308; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5309; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5310; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5311; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5312; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5313; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5314; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5315; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5316; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5317; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5318; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5319; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5320; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5321; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5322; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5323; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5324; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5325; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5326; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5327; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5328; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5329; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5330; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5331; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5332; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5333; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5334; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5335; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5336; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5337; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5338; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5339; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5340; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5341; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5342; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5343; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5344; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5345; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5346; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5347; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5348; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5349; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5350; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5351; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5352; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5353; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5354; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5355; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5356; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5357; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5358; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5359; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5360; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5361; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5362; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5363; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5364; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5365; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5366; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5367; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5368; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5369; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5370; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5371; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5372; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5373; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5374; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5375; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5376; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5377; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5378; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5379; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5380; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5381; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5382; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5383; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5384; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5385; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5386; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5387; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5388; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5389; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5390; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5391; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5392; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5393; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5394; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5395; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5396; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5397; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5398; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5399; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5400; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5401; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5402; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5403; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5404; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5405; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5406; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5407; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5408; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5409; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5410; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5411; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5412; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5413; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5414; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5415; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5416; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5417; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5418; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5419; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5420; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5421; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5422; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5423; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5424; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5425; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5426; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5427; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5428; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5429; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5430; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5431; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5432; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5433; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5434; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5435; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5436; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5437; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5438; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5439; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5440; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5441; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5442; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5443; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5444; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5445; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5446; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5447; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5448; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5449; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5450; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5451; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5452; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5453; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5454; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5455; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5456; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5457; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5458; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5459; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5460; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5461; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5462; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5463; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5464; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5465; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5466; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5467; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5468; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5469; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5470; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5471; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5472; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5473; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5474; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5475; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5476; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5477; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5478; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5479; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5480; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5481; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5482; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5483; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5484; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5485; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5486; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5487; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5488; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5489; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5490; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5491; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5492; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5493; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5494; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5495; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5496; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5497; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5498; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5499; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5500; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5501; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5502; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5503; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5504; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5505; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5506; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5507; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5508; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5509; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5510; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5511; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5512; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5513; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5514; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5515; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5516; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5517; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5518; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5519; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5520; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5521; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5522; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5523; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5524; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5525; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5526; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5527; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5528; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5529; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5530; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5531; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5532; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5533; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5534; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5535; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5536; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5537; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5538; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5539; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5540; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5541; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5542; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5543; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5544; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5545; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5546; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5547; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5548; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5549; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5550; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5551; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5552; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5553; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5554; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5555; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5556; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5557; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5558; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5559; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5560; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5561; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5562; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5563; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5564; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5565; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5566; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5567; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5568; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5569; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5570; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5571; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5572; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5573; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5574; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5575; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5576; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5577; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5578; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5579; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5580; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5581; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5582; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5583; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5584; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5585; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5586; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5587; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5588; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5589; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5590; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5591; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5592; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5593; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5594; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5595; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5596; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5597; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5598; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5599; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5600; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5601; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5602; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5603; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5604; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5605; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5606; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5607; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5608; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5609; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5610; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5611; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5612; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5613; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5614; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5615; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5616; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5617; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5618; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5619; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5620; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5621; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5622; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5623; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5624; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5625; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5626; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5627; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5628; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5629; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5630; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5631; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5632; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5633; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5634; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5635; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5636; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5637; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5638; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5639; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5640; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5641; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5642; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5643; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5644; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5645; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5646; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5647; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5648; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5649; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5650; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5651; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5652; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5653; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5654; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5655; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5656; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5657; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5658; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5659; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5660; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5661; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5662; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5663; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5664; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5665; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5666; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5667; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5668; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5669; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5670; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5671; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5672; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5673; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5674; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5675; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5676; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5677; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5678; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5679; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5680; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5681; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5682; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5683; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5684; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5685; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5686; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5687; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5688; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5689; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5690; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5691; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5692; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5693; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5694; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5695; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5696; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5697; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5698; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5699; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5700; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5701; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5702; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5703; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5704; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5705; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5706; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5707; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5708; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5709; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5710; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5711; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5712; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5713; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5714; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5715; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5716; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5717; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5718; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5719; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5720; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5721; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5722; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5723; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5724; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5725; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5726; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5727; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5728; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5729; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5730; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5731; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5732; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5733; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5734; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5735; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5736; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5737; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5738; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5739; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5740; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5741; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5742; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5743; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5744; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5745; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5746; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5747; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5748; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5749; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5750; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5751; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5752; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5753; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5754; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5755; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5756; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5757; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5758; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5759; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5760; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5761; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5762; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5763; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5764; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5765; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5766; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5767; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5768; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5769; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5770; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5771; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5772; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5773; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5774; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5775; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5776; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5777; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5778; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5779; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5780; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5781; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5782; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5783; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5784; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5785; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5786; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5787; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5788; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5789; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5790; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5791; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5792; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5793; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5794; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5795; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5796; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5797; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5798; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5799; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5800; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5801; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5802; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5803; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5804; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5805; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5806; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5807; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5808; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5809; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5810; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5811; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5812; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5813; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5814; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5815; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5816; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5817; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5818; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5819; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5820; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5821; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5822; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5823; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5824; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5825; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5826; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5827; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5828; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5829; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5830; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5831; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5832; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5833; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5834; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5835; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5836; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5837; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5838; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5839; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5840; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5841; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5842; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5843; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5844; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5845; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5846; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5847; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5848; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5849; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5850; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5851; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5852; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5853; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5854; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5855; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5856; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5857; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5858; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5859; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5860; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5861; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5862; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5863; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5864; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5865; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5866; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5867; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5868; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5869; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5870; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5871; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5872; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5873; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5874; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5875; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5876; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5877; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5878; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5879; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5880; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5881; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5882; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5883; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5884; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5885; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5886; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5887; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5888; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5889; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5890; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5891; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5892; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5893; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5894; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5895; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5896; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5897; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5898; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5899; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5900; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5901; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5902; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5903; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5904; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5905; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5906; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5907; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5908; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5909; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5910; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5911; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5912; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5913; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5914; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5915; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5916; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5917; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5918; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5919; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5920; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5921; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5922; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5923; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5924; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5925; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5926; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5927; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5928; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5929; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5930; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5931; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5932; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5933; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5934; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5935; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5936; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5937; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5938; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5939; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5940; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5941; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5942; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5943; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5944; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5945; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5946; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5947; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5948; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5949; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5950; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5951; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5952; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5953; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5954; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5955; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5956; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5957; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5958; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5959; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5960; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5961; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5962; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5963; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5964; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5965; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5966; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5967; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5968; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5969; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5970; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5971; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5972; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5973; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5974; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5975; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5976; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5977; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5978; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5979; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5980; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5981; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5982; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5983; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5984; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5985; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5986; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5987; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5988; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5989; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5990; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5991; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5992; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5993; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5994; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5995; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5996; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5997; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5998; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_5999; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_6000; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_6001; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_6002; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_6003; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_6004; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_6005; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_6006; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_6007; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_6008; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_6009; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_6010; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_6011; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_6012; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_6013; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_6014; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_6015; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_6016; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_6017; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_6018; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_6019; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_6020; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_6021; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_6022; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_6023; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_6024; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_6025; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_6026; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_6027; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_6028; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_6029; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_6030; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_6031; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_6032; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_6033; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_6034; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_6035; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_6036; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_6037; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_6038; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_6039; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_6040; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_6041; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_6042; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_6043; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_6044; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_6045; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_6046; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_6047; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_6048; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_6049; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_6050; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_6051; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_6052; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_6053; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_6054; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_6055; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_6056; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_6057; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_6058; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_6059; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_6060; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_6061; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_6062; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_6063; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_6064; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_6065; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_6066; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_6067; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_6068; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_6069; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_6070; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_6071; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_6072; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_6073; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_6074; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_6075; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_6076; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_6077; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_6078; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_6079; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_6080; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_6081; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_6082; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_6083; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_6084; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_6085; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_6086; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_6087; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_6088; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_6089; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_6090; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_6091; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_6092; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_6093; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_6094; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_6095; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_6096; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_6097; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_6098; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_6099; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_6100; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_6101; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_6102; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_6103; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_6104; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_6105; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_6106; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_6107; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_6108; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_6109; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_6110; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_6111; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_6112; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_6113; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_6114; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_6115; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_6116; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_6117; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_6118; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_6119; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_6120; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_6121; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_6122; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_6123; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_6124; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_6125; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_6126; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_6127; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_6128; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_6129; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_6130; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_6131; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_6132; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_6133; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_6134; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_6135; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_6136; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_6137; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_6138; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_6139; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_6140; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_6141; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_6142; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_6143; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_6144; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_6145; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_6146; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_6147; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_6148; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_6149; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_6150; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_6151; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_6152; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_6153; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_6154; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_6155; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_6156; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_6157; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_6158; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_6159; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_6160; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_6161; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_6162; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_6163; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_6164; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_6165; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_6166; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_6167; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_6168; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_6169; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_6170; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_6171; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_6172; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_6173; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_6174; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_6175; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_6176; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_6177; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_6178; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_6179; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_6180; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_6181; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_6182; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_6183; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_6184; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_6185; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_6186; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_6187; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_6188; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_6189; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_6190; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_6191; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_6192; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_6193; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_6194; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_6195; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_6196; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_6197; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_6198; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_6199; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_6200; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_6201; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_6202; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_6203; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_6204; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_6205; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_6206; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_6207; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_6208; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_6209; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_6210; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_6211; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_6212; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_6213; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_6214; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_6215; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_6216; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_6217; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_6218; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_6219; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_6220; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_6221; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_6222; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_6223; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_6224; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_6225; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_6226; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_6227; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_6228; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_6229; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_6230; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_6231; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_6232; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_6233; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_6234; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_6235; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_6236; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_6237; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_6238; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_6239; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_6240; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_6241; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_6242; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_6243; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_6244; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_6245; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_6246; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_6247; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_6248; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_6249; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_6250; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_6251; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_6252; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_6253; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_6254; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_6255; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_6256; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_6257; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_6258; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_6259; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_6260; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_6261; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_6262; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_6263; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_6264; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_6265; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_6266; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_6267; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_6268; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_6269; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_6270; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_6271; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_6272; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_6273; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_6274; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_6275; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_6276; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_6277; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_6278; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_6279; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_6280; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_6281; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_6282; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_6283; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_6284; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_6285; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_6286; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_6287; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_6288; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_6289; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_6290; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_6291; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_6292; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_6293; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_6294; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_6295; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_6296; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_6297; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_6298; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_6299; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_6300; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_6301; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_6302; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_6303; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_6304; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_6305; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_6306; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_6307; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_6308; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_6309; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_6310; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_6311; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_6312; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_6313; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_6314; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_6315; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_6316; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_6317; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_6318; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_6319; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_6320; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_6321; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_6322; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_6323; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_6324; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_6325; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_6326; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_6327; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_6328; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_6329; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_6330; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_6331; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_6332; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_6333; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_6334; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_6335; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_6336; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_6337; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_6338; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_6339; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_6340; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_6341; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_6342; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_6343; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_6344; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_6345; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_6346; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_6347; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_6348; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_6349; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_6350; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_6351; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_6352; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_6353; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_6354; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_6355; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_6356; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_6357; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_6358; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_6359; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_6360; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_6361; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_6362; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_6363; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_6364; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_6365; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_6366; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_6367; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_6368; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_6369; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_6370; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_6371; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_6372; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_6373; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_6374; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_6375; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_6376; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_6377; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_6378; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_6379; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_6380; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_6381; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_6382; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_6383; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_6384; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_6385; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_6386; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_6387; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_6388; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_6389; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_6390; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_6391; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_6392; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_6393; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_6394; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_6395; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_6396; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_6397; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_6398; // @[ChiselImProc.scala 188:26]
  reg [7:0] lineBuffer_6399; // @[ChiselImProc.scala 188:26]
  reg [7:0] windowBuffer_0; // @[ChiselImProc.scala 189:28]
  reg [7:0] windowBuffer_1; // @[ChiselImProc.scala 189:28]
  reg [7:0] windowBuffer_2; // @[ChiselImProc.scala 189:28]
  reg [7:0] windowBuffer_3; // @[ChiselImProc.scala 189:28]
  reg [7:0] windowBuffer_4; // @[ChiselImProc.scala 189:28]
  reg [7:0] windowBuffer_5; // @[ChiselImProc.scala 189:28]
  reg [7:0] windowBuffer_6; // @[ChiselImProc.scala 189:28]
  reg [7:0] windowBuffer_7; // @[ChiselImProc.scala 189:28]
  reg [7:0] windowBuffer_8; // @[ChiselImProc.scala 189:28]
  reg [7:0] windowBuffer_9; // @[ChiselImProc.scala 189:28]
  reg [7:0] windowBuffer_10; // @[ChiselImProc.scala 189:28]
  reg [7:0] windowBuffer_11; // @[ChiselImProc.scala 189:28]
  reg [7:0] windowBuffer_12; // @[ChiselImProc.scala 189:28]
  reg [7:0] windowBuffer_13; // @[ChiselImProc.scala 189:28]
  reg [7:0] windowBuffer_14; // @[ChiselImProc.scala 189:28]
  reg [7:0] windowBuffer_15; // @[ChiselImProc.scala 189:28]
  reg [7:0] windowBuffer_16; // @[ChiselImProc.scala 189:28]
  reg [7:0] windowBuffer_17; // @[ChiselImProc.scala 189:28]
  reg [7:0] windowBuffer_18; // @[ChiselImProc.scala 189:28]
  reg [7:0] windowBuffer_19; // @[ChiselImProc.scala 189:28]
  reg [7:0] windowBuffer_20; // @[ChiselImProc.scala 189:28]
  reg [7:0] windowBuffer_21; // @[ChiselImProc.scala 189:28]
  reg [7:0] windowBuffer_22; // @[ChiselImProc.scala 189:28]
  reg [7:0] windowBuffer_23; // @[ChiselImProc.scala 189:28]
  reg [7:0] windowBuffer_24; // @[ChiselImProc.scala 189:28]
  wire  sel = _T_16 & io_deq_ready; // @[ChiselImProc.scala 192:47]
  MulAdd MulAdd ( // @[ChiselImProc.scala 206:29]
    .io_b_0(MulAdd_io_b_0),
    .io_b_1(MulAdd_io_b_1),
    .io_b_2(MulAdd_io_b_2),
    .io_b_3(MulAdd_io_b_3),
    .io_b_4(MulAdd_io_b_4),
    .io_b_5(MulAdd_io_b_5),
    .io_b_6(MulAdd_io_b_6),
    .io_b_7(MulAdd_io_b_7),
    .io_b_8(MulAdd_io_b_8),
    .io_b_9(MulAdd_io_b_9),
    .io_b_10(MulAdd_io_b_10),
    .io_b_11(MulAdd_io_b_11),
    .io_b_12(MulAdd_io_b_12),
    .io_b_13(MulAdd_io_b_13),
    .io_b_14(MulAdd_io_b_14),
    .io_b_15(MulAdd_io_b_15),
    .io_b_16(MulAdd_io_b_16),
    .io_b_17(MulAdd_io_b_17),
    .io_b_18(MulAdd_io_b_18),
    .io_b_19(MulAdd_io_b_19),
    .io_b_20(MulAdd_io_b_20),
    .io_b_21(MulAdd_io_b_21),
    .io_b_22(MulAdd_io_b_22),
    .io_b_23(MulAdd_io_b_23),
    .io_b_24(MulAdd_io_b_24),
    .io_output(MulAdd_io_output)
  );
  assign io_enq_ready = _T_11 | _T_12; // @[ChiselImProc.scala 110:22]
  assign io_deq_valid = _T_10 | _T_15; // @[ChiselImProc.scala 111:22]
  assign io_deq_bits = MulAdd_io_output[15:8]; // @[ChiselImProc.scala 211:17]
  assign io_deq_user = userReg; // @[ChiselImProc.scala 138:17 ChiselImProc.scala 108:21]
  assign io_deq_last = lastReg; // @[ChiselImProc.scala 137:17 ChiselImProc.scala 107:21]
  assign MulAdd_io_b_0 = windowBuffer_0; // @[ChiselImProc.scala 209:13]
  assign MulAdd_io_b_1 = windowBuffer_1; // @[ChiselImProc.scala 209:13]
  assign MulAdd_io_b_2 = windowBuffer_2; // @[ChiselImProc.scala 209:13]
  assign MulAdd_io_b_3 = windowBuffer_3; // @[ChiselImProc.scala 209:13]
  assign MulAdd_io_b_4 = windowBuffer_4; // @[ChiselImProc.scala 209:13]
  assign MulAdd_io_b_5 = windowBuffer_5; // @[ChiselImProc.scala 209:13]
  assign MulAdd_io_b_6 = windowBuffer_6; // @[ChiselImProc.scala 209:13]
  assign MulAdd_io_b_7 = windowBuffer_7; // @[ChiselImProc.scala 209:13]
  assign MulAdd_io_b_8 = windowBuffer_8; // @[ChiselImProc.scala 209:13]
  assign MulAdd_io_b_9 = windowBuffer_9; // @[ChiselImProc.scala 209:13]
  assign MulAdd_io_b_10 = windowBuffer_10; // @[ChiselImProc.scala 209:13]
  assign MulAdd_io_b_11 = windowBuffer_11; // @[ChiselImProc.scala 209:13]
  assign MulAdd_io_b_12 = windowBuffer_12; // @[ChiselImProc.scala 209:13]
  assign MulAdd_io_b_13 = windowBuffer_13; // @[ChiselImProc.scala 209:13]
  assign MulAdd_io_b_14 = windowBuffer_14; // @[ChiselImProc.scala 209:13]
  assign MulAdd_io_b_15 = windowBuffer_15; // @[ChiselImProc.scala 209:13]
  assign MulAdd_io_b_16 = windowBuffer_16; // @[ChiselImProc.scala 209:13]
  assign MulAdd_io_b_17 = windowBuffer_17; // @[ChiselImProc.scala 209:13]
  assign MulAdd_io_b_18 = windowBuffer_18; // @[ChiselImProc.scala 209:13]
  assign MulAdd_io_b_19 = windowBuffer_19; // @[ChiselImProc.scala 209:13]
  assign MulAdd_io_b_20 = windowBuffer_20; // @[ChiselImProc.scala 209:13]
  assign MulAdd_io_b_21 = windowBuffer_21; // @[ChiselImProc.scala 209:13]
  assign MulAdd_io_b_22 = windowBuffer_22; // @[ChiselImProc.scala 209:13]
  assign MulAdd_io_b_23 = windowBuffer_23; // @[ChiselImProc.scala 209:13]
  assign MulAdd_io_b_24 = windowBuffer_24; // @[ChiselImProc.scala 209:13]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  stateReg = _RAND_0[1:0];
  _RAND_1 = {1{`RANDOM}};
  dataReg = _RAND_1[7:0];
  _RAND_2 = {1{`RANDOM}};
  shadowReg = _RAND_2[7:0];
  _RAND_3 = {1{`RANDOM}};
  userReg = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  shadowUserReg = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  lastReg = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  shadowLastReg = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  lineBuffer_0 = _RAND_7[7:0];
  _RAND_8 = {1{`RANDOM}};
  lineBuffer_1 = _RAND_8[7:0];
  _RAND_9 = {1{`RANDOM}};
  lineBuffer_2 = _RAND_9[7:0];
  _RAND_10 = {1{`RANDOM}};
  lineBuffer_3 = _RAND_10[7:0];
  _RAND_11 = {1{`RANDOM}};
  lineBuffer_4 = _RAND_11[7:0];
  _RAND_12 = {1{`RANDOM}};
  lineBuffer_5 = _RAND_12[7:0];
  _RAND_13 = {1{`RANDOM}};
  lineBuffer_6 = _RAND_13[7:0];
  _RAND_14 = {1{`RANDOM}};
  lineBuffer_7 = _RAND_14[7:0];
  _RAND_15 = {1{`RANDOM}};
  lineBuffer_8 = _RAND_15[7:0];
  _RAND_16 = {1{`RANDOM}};
  lineBuffer_9 = _RAND_16[7:0];
  _RAND_17 = {1{`RANDOM}};
  lineBuffer_10 = _RAND_17[7:0];
  _RAND_18 = {1{`RANDOM}};
  lineBuffer_11 = _RAND_18[7:0];
  _RAND_19 = {1{`RANDOM}};
  lineBuffer_12 = _RAND_19[7:0];
  _RAND_20 = {1{`RANDOM}};
  lineBuffer_13 = _RAND_20[7:0];
  _RAND_21 = {1{`RANDOM}};
  lineBuffer_14 = _RAND_21[7:0];
  _RAND_22 = {1{`RANDOM}};
  lineBuffer_15 = _RAND_22[7:0];
  _RAND_23 = {1{`RANDOM}};
  lineBuffer_16 = _RAND_23[7:0];
  _RAND_24 = {1{`RANDOM}};
  lineBuffer_17 = _RAND_24[7:0];
  _RAND_25 = {1{`RANDOM}};
  lineBuffer_18 = _RAND_25[7:0];
  _RAND_26 = {1{`RANDOM}};
  lineBuffer_19 = _RAND_26[7:0];
  _RAND_27 = {1{`RANDOM}};
  lineBuffer_20 = _RAND_27[7:0];
  _RAND_28 = {1{`RANDOM}};
  lineBuffer_21 = _RAND_28[7:0];
  _RAND_29 = {1{`RANDOM}};
  lineBuffer_22 = _RAND_29[7:0];
  _RAND_30 = {1{`RANDOM}};
  lineBuffer_23 = _RAND_30[7:0];
  _RAND_31 = {1{`RANDOM}};
  lineBuffer_24 = _RAND_31[7:0];
  _RAND_32 = {1{`RANDOM}};
  lineBuffer_25 = _RAND_32[7:0];
  _RAND_33 = {1{`RANDOM}};
  lineBuffer_26 = _RAND_33[7:0];
  _RAND_34 = {1{`RANDOM}};
  lineBuffer_27 = _RAND_34[7:0];
  _RAND_35 = {1{`RANDOM}};
  lineBuffer_28 = _RAND_35[7:0];
  _RAND_36 = {1{`RANDOM}};
  lineBuffer_29 = _RAND_36[7:0];
  _RAND_37 = {1{`RANDOM}};
  lineBuffer_30 = _RAND_37[7:0];
  _RAND_38 = {1{`RANDOM}};
  lineBuffer_31 = _RAND_38[7:0];
  _RAND_39 = {1{`RANDOM}};
  lineBuffer_32 = _RAND_39[7:0];
  _RAND_40 = {1{`RANDOM}};
  lineBuffer_33 = _RAND_40[7:0];
  _RAND_41 = {1{`RANDOM}};
  lineBuffer_34 = _RAND_41[7:0];
  _RAND_42 = {1{`RANDOM}};
  lineBuffer_35 = _RAND_42[7:0];
  _RAND_43 = {1{`RANDOM}};
  lineBuffer_36 = _RAND_43[7:0];
  _RAND_44 = {1{`RANDOM}};
  lineBuffer_37 = _RAND_44[7:0];
  _RAND_45 = {1{`RANDOM}};
  lineBuffer_38 = _RAND_45[7:0];
  _RAND_46 = {1{`RANDOM}};
  lineBuffer_39 = _RAND_46[7:0];
  _RAND_47 = {1{`RANDOM}};
  lineBuffer_40 = _RAND_47[7:0];
  _RAND_48 = {1{`RANDOM}};
  lineBuffer_41 = _RAND_48[7:0];
  _RAND_49 = {1{`RANDOM}};
  lineBuffer_42 = _RAND_49[7:0];
  _RAND_50 = {1{`RANDOM}};
  lineBuffer_43 = _RAND_50[7:0];
  _RAND_51 = {1{`RANDOM}};
  lineBuffer_44 = _RAND_51[7:0];
  _RAND_52 = {1{`RANDOM}};
  lineBuffer_45 = _RAND_52[7:0];
  _RAND_53 = {1{`RANDOM}};
  lineBuffer_46 = _RAND_53[7:0];
  _RAND_54 = {1{`RANDOM}};
  lineBuffer_47 = _RAND_54[7:0];
  _RAND_55 = {1{`RANDOM}};
  lineBuffer_48 = _RAND_55[7:0];
  _RAND_56 = {1{`RANDOM}};
  lineBuffer_49 = _RAND_56[7:0];
  _RAND_57 = {1{`RANDOM}};
  lineBuffer_50 = _RAND_57[7:0];
  _RAND_58 = {1{`RANDOM}};
  lineBuffer_51 = _RAND_58[7:0];
  _RAND_59 = {1{`RANDOM}};
  lineBuffer_52 = _RAND_59[7:0];
  _RAND_60 = {1{`RANDOM}};
  lineBuffer_53 = _RAND_60[7:0];
  _RAND_61 = {1{`RANDOM}};
  lineBuffer_54 = _RAND_61[7:0];
  _RAND_62 = {1{`RANDOM}};
  lineBuffer_55 = _RAND_62[7:0];
  _RAND_63 = {1{`RANDOM}};
  lineBuffer_56 = _RAND_63[7:0];
  _RAND_64 = {1{`RANDOM}};
  lineBuffer_57 = _RAND_64[7:0];
  _RAND_65 = {1{`RANDOM}};
  lineBuffer_58 = _RAND_65[7:0];
  _RAND_66 = {1{`RANDOM}};
  lineBuffer_59 = _RAND_66[7:0];
  _RAND_67 = {1{`RANDOM}};
  lineBuffer_60 = _RAND_67[7:0];
  _RAND_68 = {1{`RANDOM}};
  lineBuffer_61 = _RAND_68[7:0];
  _RAND_69 = {1{`RANDOM}};
  lineBuffer_62 = _RAND_69[7:0];
  _RAND_70 = {1{`RANDOM}};
  lineBuffer_63 = _RAND_70[7:0];
  _RAND_71 = {1{`RANDOM}};
  lineBuffer_64 = _RAND_71[7:0];
  _RAND_72 = {1{`RANDOM}};
  lineBuffer_65 = _RAND_72[7:0];
  _RAND_73 = {1{`RANDOM}};
  lineBuffer_66 = _RAND_73[7:0];
  _RAND_74 = {1{`RANDOM}};
  lineBuffer_67 = _RAND_74[7:0];
  _RAND_75 = {1{`RANDOM}};
  lineBuffer_68 = _RAND_75[7:0];
  _RAND_76 = {1{`RANDOM}};
  lineBuffer_69 = _RAND_76[7:0];
  _RAND_77 = {1{`RANDOM}};
  lineBuffer_70 = _RAND_77[7:0];
  _RAND_78 = {1{`RANDOM}};
  lineBuffer_71 = _RAND_78[7:0];
  _RAND_79 = {1{`RANDOM}};
  lineBuffer_72 = _RAND_79[7:0];
  _RAND_80 = {1{`RANDOM}};
  lineBuffer_73 = _RAND_80[7:0];
  _RAND_81 = {1{`RANDOM}};
  lineBuffer_74 = _RAND_81[7:0];
  _RAND_82 = {1{`RANDOM}};
  lineBuffer_75 = _RAND_82[7:0];
  _RAND_83 = {1{`RANDOM}};
  lineBuffer_76 = _RAND_83[7:0];
  _RAND_84 = {1{`RANDOM}};
  lineBuffer_77 = _RAND_84[7:0];
  _RAND_85 = {1{`RANDOM}};
  lineBuffer_78 = _RAND_85[7:0];
  _RAND_86 = {1{`RANDOM}};
  lineBuffer_79 = _RAND_86[7:0];
  _RAND_87 = {1{`RANDOM}};
  lineBuffer_80 = _RAND_87[7:0];
  _RAND_88 = {1{`RANDOM}};
  lineBuffer_81 = _RAND_88[7:0];
  _RAND_89 = {1{`RANDOM}};
  lineBuffer_82 = _RAND_89[7:0];
  _RAND_90 = {1{`RANDOM}};
  lineBuffer_83 = _RAND_90[7:0];
  _RAND_91 = {1{`RANDOM}};
  lineBuffer_84 = _RAND_91[7:0];
  _RAND_92 = {1{`RANDOM}};
  lineBuffer_85 = _RAND_92[7:0];
  _RAND_93 = {1{`RANDOM}};
  lineBuffer_86 = _RAND_93[7:0];
  _RAND_94 = {1{`RANDOM}};
  lineBuffer_87 = _RAND_94[7:0];
  _RAND_95 = {1{`RANDOM}};
  lineBuffer_88 = _RAND_95[7:0];
  _RAND_96 = {1{`RANDOM}};
  lineBuffer_89 = _RAND_96[7:0];
  _RAND_97 = {1{`RANDOM}};
  lineBuffer_90 = _RAND_97[7:0];
  _RAND_98 = {1{`RANDOM}};
  lineBuffer_91 = _RAND_98[7:0];
  _RAND_99 = {1{`RANDOM}};
  lineBuffer_92 = _RAND_99[7:0];
  _RAND_100 = {1{`RANDOM}};
  lineBuffer_93 = _RAND_100[7:0];
  _RAND_101 = {1{`RANDOM}};
  lineBuffer_94 = _RAND_101[7:0];
  _RAND_102 = {1{`RANDOM}};
  lineBuffer_95 = _RAND_102[7:0];
  _RAND_103 = {1{`RANDOM}};
  lineBuffer_96 = _RAND_103[7:0];
  _RAND_104 = {1{`RANDOM}};
  lineBuffer_97 = _RAND_104[7:0];
  _RAND_105 = {1{`RANDOM}};
  lineBuffer_98 = _RAND_105[7:0];
  _RAND_106 = {1{`RANDOM}};
  lineBuffer_99 = _RAND_106[7:0];
  _RAND_107 = {1{`RANDOM}};
  lineBuffer_100 = _RAND_107[7:0];
  _RAND_108 = {1{`RANDOM}};
  lineBuffer_101 = _RAND_108[7:0];
  _RAND_109 = {1{`RANDOM}};
  lineBuffer_102 = _RAND_109[7:0];
  _RAND_110 = {1{`RANDOM}};
  lineBuffer_103 = _RAND_110[7:0];
  _RAND_111 = {1{`RANDOM}};
  lineBuffer_104 = _RAND_111[7:0];
  _RAND_112 = {1{`RANDOM}};
  lineBuffer_105 = _RAND_112[7:0];
  _RAND_113 = {1{`RANDOM}};
  lineBuffer_106 = _RAND_113[7:0];
  _RAND_114 = {1{`RANDOM}};
  lineBuffer_107 = _RAND_114[7:0];
  _RAND_115 = {1{`RANDOM}};
  lineBuffer_108 = _RAND_115[7:0];
  _RAND_116 = {1{`RANDOM}};
  lineBuffer_109 = _RAND_116[7:0];
  _RAND_117 = {1{`RANDOM}};
  lineBuffer_110 = _RAND_117[7:0];
  _RAND_118 = {1{`RANDOM}};
  lineBuffer_111 = _RAND_118[7:0];
  _RAND_119 = {1{`RANDOM}};
  lineBuffer_112 = _RAND_119[7:0];
  _RAND_120 = {1{`RANDOM}};
  lineBuffer_113 = _RAND_120[7:0];
  _RAND_121 = {1{`RANDOM}};
  lineBuffer_114 = _RAND_121[7:0];
  _RAND_122 = {1{`RANDOM}};
  lineBuffer_115 = _RAND_122[7:0];
  _RAND_123 = {1{`RANDOM}};
  lineBuffer_116 = _RAND_123[7:0];
  _RAND_124 = {1{`RANDOM}};
  lineBuffer_117 = _RAND_124[7:0];
  _RAND_125 = {1{`RANDOM}};
  lineBuffer_118 = _RAND_125[7:0];
  _RAND_126 = {1{`RANDOM}};
  lineBuffer_119 = _RAND_126[7:0];
  _RAND_127 = {1{`RANDOM}};
  lineBuffer_120 = _RAND_127[7:0];
  _RAND_128 = {1{`RANDOM}};
  lineBuffer_121 = _RAND_128[7:0];
  _RAND_129 = {1{`RANDOM}};
  lineBuffer_122 = _RAND_129[7:0];
  _RAND_130 = {1{`RANDOM}};
  lineBuffer_123 = _RAND_130[7:0];
  _RAND_131 = {1{`RANDOM}};
  lineBuffer_124 = _RAND_131[7:0];
  _RAND_132 = {1{`RANDOM}};
  lineBuffer_125 = _RAND_132[7:0];
  _RAND_133 = {1{`RANDOM}};
  lineBuffer_126 = _RAND_133[7:0];
  _RAND_134 = {1{`RANDOM}};
  lineBuffer_127 = _RAND_134[7:0];
  _RAND_135 = {1{`RANDOM}};
  lineBuffer_128 = _RAND_135[7:0];
  _RAND_136 = {1{`RANDOM}};
  lineBuffer_129 = _RAND_136[7:0];
  _RAND_137 = {1{`RANDOM}};
  lineBuffer_130 = _RAND_137[7:0];
  _RAND_138 = {1{`RANDOM}};
  lineBuffer_131 = _RAND_138[7:0];
  _RAND_139 = {1{`RANDOM}};
  lineBuffer_132 = _RAND_139[7:0];
  _RAND_140 = {1{`RANDOM}};
  lineBuffer_133 = _RAND_140[7:0];
  _RAND_141 = {1{`RANDOM}};
  lineBuffer_134 = _RAND_141[7:0];
  _RAND_142 = {1{`RANDOM}};
  lineBuffer_135 = _RAND_142[7:0];
  _RAND_143 = {1{`RANDOM}};
  lineBuffer_136 = _RAND_143[7:0];
  _RAND_144 = {1{`RANDOM}};
  lineBuffer_137 = _RAND_144[7:0];
  _RAND_145 = {1{`RANDOM}};
  lineBuffer_138 = _RAND_145[7:0];
  _RAND_146 = {1{`RANDOM}};
  lineBuffer_139 = _RAND_146[7:0];
  _RAND_147 = {1{`RANDOM}};
  lineBuffer_140 = _RAND_147[7:0];
  _RAND_148 = {1{`RANDOM}};
  lineBuffer_141 = _RAND_148[7:0];
  _RAND_149 = {1{`RANDOM}};
  lineBuffer_142 = _RAND_149[7:0];
  _RAND_150 = {1{`RANDOM}};
  lineBuffer_143 = _RAND_150[7:0];
  _RAND_151 = {1{`RANDOM}};
  lineBuffer_144 = _RAND_151[7:0];
  _RAND_152 = {1{`RANDOM}};
  lineBuffer_145 = _RAND_152[7:0];
  _RAND_153 = {1{`RANDOM}};
  lineBuffer_146 = _RAND_153[7:0];
  _RAND_154 = {1{`RANDOM}};
  lineBuffer_147 = _RAND_154[7:0];
  _RAND_155 = {1{`RANDOM}};
  lineBuffer_148 = _RAND_155[7:0];
  _RAND_156 = {1{`RANDOM}};
  lineBuffer_149 = _RAND_156[7:0];
  _RAND_157 = {1{`RANDOM}};
  lineBuffer_150 = _RAND_157[7:0];
  _RAND_158 = {1{`RANDOM}};
  lineBuffer_151 = _RAND_158[7:0];
  _RAND_159 = {1{`RANDOM}};
  lineBuffer_152 = _RAND_159[7:0];
  _RAND_160 = {1{`RANDOM}};
  lineBuffer_153 = _RAND_160[7:0];
  _RAND_161 = {1{`RANDOM}};
  lineBuffer_154 = _RAND_161[7:0];
  _RAND_162 = {1{`RANDOM}};
  lineBuffer_155 = _RAND_162[7:0];
  _RAND_163 = {1{`RANDOM}};
  lineBuffer_156 = _RAND_163[7:0];
  _RAND_164 = {1{`RANDOM}};
  lineBuffer_157 = _RAND_164[7:0];
  _RAND_165 = {1{`RANDOM}};
  lineBuffer_158 = _RAND_165[7:0];
  _RAND_166 = {1{`RANDOM}};
  lineBuffer_159 = _RAND_166[7:0];
  _RAND_167 = {1{`RANDOM}};
  lineBuffer_160 = _RAND_167[7:0];
  _RAND_168 = {1{`RANDOM}};
  lineBuffer_161 = _RAND_168[7:0];
  _RAND_169 = {1{`RANDOM}};
  lineBuffer_162 = _RAND_169[7:0];
  _RAND_170 = {1{`RANDOM}};
  lineBuffer_163 = _RAND_170[7:0];
  _RAND_171 = {1{`RANDOM}};
  lineBuffer_164 = _RAND_171[7:0];
  _RAND_172 = {1{`RANDOM}};
  lineBuffer_165 = _RAND_172[7:0];
  _RAND_173 = {1{`RANDOM}};
  lineBuffer_166 = _RAND_173[7:0];
  _RAND_174 = {1{`RANDOM}};
  lineBuffer_167 = _RAND_174[7:0];
  _RAND_175 = {1{`RANDOM}};
  lineBuffer_168 = _RAND_175[7:0];
  _RAND_176 = {1{`RANDOM}};
  lineBuffer_169 = _RAND_176[7:0];
  _RAND_177 = {1{`RANDOM}};
  lineBuffer_170 = _RAND_177[7:0];
  _RAND_178 = {1{`RANDOM}};
  lineBuffer_171 = _RAND_178[7:0];
  _RAND_179 = {1{`RANDOM}};
  lineBuffer_172 = _RAND_179[7:0];
  _RAND_180 = {1{`RANDOM}};
  lineBuffer_173 = _RAND_180[7:0];
  _RAND_181 = {1{`RANDOM}};
  lineBuffer_174 = _RAND_181[7:0];
  _RAND_182 = {1{`RANDOM}};
  lineBuffer_175 = _RAND_182[7:0];
  _RAND_183 = {1{`RANDOM}};
  lineBuffer_176 = _RAND_183[7:0];
  _RAND_184 = {1{`RANDOM}};
  lineBuffer_177 = _RAND_184[7:0];
  _RAND_185 = {1{`RANDOM}};
  lineBuffer_178 = _RAND_185[7:0];
  _RAND_186 = {1{`RANDOM}};
  lineBuffer_179 = _RAND_186[7:0];
  _RAND_187 = {1{`RANDOM}};
  lineBuffer_180 = _RAND_187[7:0];
  _RAND_188 = {1{`RANDOM}};
  lineBuffer_181 = _RAND_188[7:0];
  _RAND_189 = {1{`RANDOM}};
  lineBuffer_182 = _RAND_189[7:0];
  _RAND_190 = {1{`RANDOM}};
  lineBuffer_183 = _RAND_190[7:0];
  _RAND_191 = {1{`RANDOM}};
  lineBuffer_184 = _RAND_191[7:0];
  _RAND_192 = {1{`RANDOM}};
  lineBuffer_185 = _RAND_192[7:0];
  _RAND_193 = {1{`RANDOM}};
  lineBuffer_186 = _RAND_193[7:0];
  _RAND_194 = {1{`RANDOM}};
  lineBuffer_187 = _RAND_194[7:0];
  _RAND_195 = {1{`RANDOM}};
  lineBuffer_188 = _RAND_195[7:0];
  _RAND_196 = {1{`RANDOM}};
  lineBuffer_189 = _RAND_196[7:0];
  _RAND_197 = {1{`RANDOM}};
  lineBuffer_190 = _RAND_197[7:0];
  _RAND_198 = {1{`RANDOM}};
  lineBuffer_191 = _RAND_198[7:0];
  _RAND_199 = {1{`RANDOM}};
  lineBuffer_192 = _RAND_199[7:0];
  _RAND_200 = {1{`RANDOM}};
  lineBuffer_193 = _RAND_200[7:0];
  _RAND_201 = {1{`RANDOM}};
  lineBuffer_194 = _RAND_201[7:0];
  _RAND_202 = {1{`RANDOM}};
  lineBuffer_195 = _RAND_202[7:0];
  _RAND_203 = {1{`RANDOM}};
  lineBuffer_196 = _RAND_203[7:0];
  _RAND_204 = {1{`RANDOM}};
  lineBuffer_197 = _RAND_204[7:0];
  _RAND_205 = {1{`RANDOM}};
  lineBuffer_198 = _RAND_205[7:0];
  _RAND_206 = {1{`RANDOM}};
  lineBuffer_199 = _RAND_206[7:0];
  _RAND_207 = {1{`RANDOM}};
  lineBuffer_200 = _RAND_207[7:0];
  _RAND_208 = {1{`RANDOM}};
  lineBuffer_201 = _RAND_208[7:0];
  _RAND_209 = {1{`RANDOM}};
  lineBuffer_202 = _RAND_209[7:0];
  _RAND_210 = {1{`RANDOM}};
  lineBuffer_203 = _RAND_210[7:0];
  _RAND_211 = {1{`RANDOM}};
  lineBuffer_204 = _RAND_211[7:0];
  _RAND_212 = {1{`RANDOM}};
  lineBuffer_205 = _RAND_212[7:0];
  _RAND_213 = {1{`RANDOM}};
  lineBuffer_206 = _RAND_213[7:0];
  _RAND_214 = {1{`RANDOM}};
  lineBuffer_207 = _RAND_214[7:0];
  _RAND_215 = {1{`RANDOM}};
  lineBuffer_208 = _RAND_215[7:0];
  _RAND_216 = {1{`RANDOM}};
  lineBuffer_209 = _RAND_216[7:0];
  _RAND_217 = {1{`RANDOM}};
  lineBuffer_210 = _RAND_217[7:0];
  _RAND_218 = {1{`RANDOM}};
  lineBuffer_211 = _RAND_218[7:0];
  _RAND_219 = {1{`RANDOM}};
  lineBuffer_212 = _RAND_219[7:0];
  _RAND_220 = {1{`RANDOM}};
  lineBuffer_213 = _RAND_220[7:0];
  _RAND_221 = {1{`RANDOM}};
  lineBuffer_214 = _RAND_221[7:0];
  _RAND_222 = {1{`RANDOM}};
  lineBuffer_215 = _RAND_222[7:0];
  _RAND_223 = {1{`RANDOM}};
  lineBuffer_216 = _RAND_223[7:0];
  _RAND_224 = {1{`RANDOM}};
  lineBuffer_217 = _RAND_224[7:0];
  _RAND_225 = {1{`RANDOM}};
  lineBuffer_218 = _RAND_225[7:0];
  _RAND_226 = {1{`RANDOM}};
  lineBuffer_219 = _RAND_226[7:0];
  _RAND_227 = {1{`RANDOM}};
  lineBuffer_220 = _RAND_227[7:0];
  _RAND_228 = {1{`RANDOM}};
  lineBuffer_221 = _RAND_228[7:0];
  _RAND_229 = {1{`RANDOM}};
  lineBuffer_222 = _RAND_229[7:0];
  _RAND_230 = {1{`RANDOM}};
  lineBuffer_223 = _RAND_230[7:0];
  _RAND_231 = {1{`RANDOM}};
  lineBuffer_224 = _RAND_231[7:0];
  _RAND_232 = {1{`RANDOM}};
  lineBuffer_225 = _RAND_232[7:0];
  _RAND_233 = {1{`RANDOM}};
  lineBuffer_226 = _RAND_233[7:0];
  _RAND_234 = {1{`RANDOM}};
  lineBuffer_227 = _RAND_234[7:0];
  _RAND_235 = {1{`RANDOM}};
  lineBuffer_228 = _RAND_235[7:0];
  _RAND_236 = {1{`RANDOM}};
  lineBuffer_229 = _RAND_236[7:0];
  _RAND_237 = {1{`RANDOM}};
  lineBuffer_230 = _RAND_237[7:0];
  _RAND_238 = {1{`RANDOM}};
  lineBuffer_231 = _RAND_238[7:0];
  _RAND_239 = {1{`RANDOM}};
  lineBuffer_232 = _RAND_239[7:0];
  _RAND_240 = {1{`RANDOM}};
  lineBuffer_233 = _RAND_240[7:0];
  _RAND_241 = {1{`RANDOM}};
  lineBuffer_234 = _RAND_241[7:0];
  _RAND_242 = {1{`RANDOM}};
  lineBuffer_235 = _RAND_242[7:0];
  _RAND_243 = {1{`RANDOM}};
  lineBuffer_236 = _RAND_243[7:0];
  _RAND_244 = {1{`RANDOM}};
  lineBuffer_237 = _RAND_244[7:0];
  _RAND_245 = {1{`RANDOM}};
  lineBuffer_238 = _RAND_245[7:0];
  _RAND_246 = {1{`RANDOM}};
  lineBuffer_239 = _RAND_246[7:0];
  _RAND_247 = {1{`RANDOM}};
  lineBuffer_240 = _RAND_247[7:0];
  _RAND_248 = {1{`RANDOM}};
  lineBuffer_241 = _RAND_248[7:0];
  _RAND_249 = {1{`RANDOM}};
  lineBuffer_242 = _RAND_249[7:0];
  _RAND_250 = {1{`RANDOM}};
  lineBuffer_243 = _RAND_250[7:0];
  _RAND_251 = {1{`RANDOM}};
  lineBuffer_244 = _RAND_251[7:0];
  _RAND_252 = {1{`RANDOM}};
  lineBuffer_245 = _RAND_252[7:0];
  _RAND_253 = {1{`RANDOM}};
  lineBuffer_246 = _RAND_253[7:0];
  _RAND_254 = {1{`RANDOM}};
  lineBuffer_247 = _RAND_254[7:0];
  _RAND_255 = {1{`RANDOM}};
  lineBuffer_248 = _RAND_255[7:0];
  _RAND_256 = {1{`RANDOM}};
  lineBuffer_249 = _RAND_256[7:0];
  _RAND_257 = {1{`RANDOM}};
  lineBuffer_250 = _RAND_257[7:0];
  _RAND_258 = {1{`RANDOM}};
  lineBuffer_251 = _RAND_258[7:0];
  _RAND_259 = {1{`RANDOM}};
  lineBuffer_252 = _RAND_259[7:0];
  _RAND_260 = {1{`RANDOM}};
  lineBuffer_253 = _RAND_260[7:0];
  _RAND_261 = {1{`RANDOM}};
  lineBuffer_254 = _RAND_261[7:0];
  _RAND_262 = {1{`RANDOM}};
  lineBuffer_255 = _RAND_262[7:0];
  _RAND_263 = {1{`RANDOM}};
  lineBuffer_256 = _RAND_263[7:0];
  _RAND_264 = {1{`RANDOM}};
  lineBuffer_257 = _RAND_264[7:0];
  _RAND_265 = {1{`RANDOM}};
  lineBuffer_258 = _RAND_265[7:0];
  _RAND_266 = {1{`RANDOM}};
  lineBuffer_259 = _RAND_266[7:0];
  _RAND_267 = {1{`RANDOM}};
  lineBuffer_260 = _RAND_267[7:0];
  _RAND_268 = {1{`RANDOM}};
  lineBuffer_261 = _RAND_268[7:0];
  _RAND_269 = {1{`RANDOM}};
  lineBuffer_262 = _RAND_269[7:0];
  _RAND_270 = {1{`RANDOM}};
  lineBuffer_263 = _RAND_270[7:0];
  _RAND_271 = {1{`RANDOM}};
  lineBuffer_264 = _RAND_271[7:0];
  _RAND_272 = {1{`RANDOM}};
  lineBuffer_265 = _RAND_272[7:0];
  _RAND_273 = {1{`RANDOM}};
  lineBuffer_266 = _RAND_273[7:0];
  _RAND_274 = {1{`RANDOM}};
  lineBuffer_267 = _RAND_274[7:0];
  _RAND_275 = {1{`RANDOM}};
  lineBuffer_268 = _RAND_275[7:0];
  _RAND_276 = {1{`RANDOM}};
  lineBuffer_269 = _RAND_276[7:0];
  _RAND_277 = {1{`RANDOM}};
  lineBuffer_270 = _RAND_277[7:0];
  _RAND_278 = {1{`RANDOM}};
  lineBuffer_271 = _RAND_278[7:0];
  _RAND_279 = {1{`RANDOM}};
  lineBuffer_272 = _RAND_279[7:0];
  _RAND_280 = {1{`RANDOM}};
  lineBuffer_273 = _RAND_280[7:0];
  _RAND_281 = {1{`RANDOM}};
  lineBuffer_274 = _RAND_281[7:0];
  _RAND_282 = {1{`RANDOM}};
  lineBuffer_275 = _RAND_282[7:0];
  _RAND_283 = {1{`RANDOM}};
  lineBuffer_276 = _RAND_283[7:0];
  _RAND_284 = {1{`RANDOM}};
  lineBuffer_277 = _RAND_284[7:0];
  _RAND_285 = {1{`RANDOM}};
  lineBuffer_278 = _RAND_285[7:0];
  _RAND_286 = {1{`RANDOM}};
  lineBuffer_279 = _RAND_286[7:0];
  _RAND_287 = {1{`RANDOM}};
  lineBuffer_280 = _RAND_287[7:0];
  _RAND_288 = {1{`RANDOM}};
  lineBuffer_281 = _RAND_288[7:0];
  _RAND_289 = {1{`RANDOM}};
  lineBuffer_282 = _RAND_289[7:0];
  _RAND_290 = {1{`RANDOM}};
  lineBuffer_283 = _RAND_290[7:0];
  _RAND_291 = {1{`RANDOM}};
  lineBuffer_284 = _RAND_291[7:0];
  _RAND_292 = {1{`RANDOM}};
  lineBuffer_285 = _RAND_292[7:0];
  _RAND_293 = {1{`RANDOM}};
  lineBuffer_286 = _RAND_293[7:0];
  _RAND_294 = {1{`RANDOM}};
  lineBuffer_287 = _RAND_294[7:0];
  _RAND_295 = {1{`RANDOM}};
  lineBuffer_288 = _RAND_295[7:0];
  _RAND_296 = {1{`RANDOM}};
  lineBuffer_289 = _RAND_296[7:0];
  _RAND_297 = {1{`RANDOM}};
  lineBuffer_290 = _RAND_297[7:0];
  _RAND_298 = {1{`RANDOM}};
  lineBuffer_291 = _RAND_298[7:0];
  _RAND_299 = {1{`RANDOM}};
  lineBuffer_292 = _RAND_299[7:0];
  _RAND_300 = {1{`RANDOM}};
  lineBuffer_293 = _RAND_300[7:0];
  _RAND_301 = {1{`RANDOM}};
  lineBuffer_294 = _RAND_301[7:0];
  _RAND_302 = {1{`RANDOM}};
  lineBuffer_295 = _RAND_302[7:0];
  _RAND_303 = {1{`RANDOM}};
  lineBuffer_296 = _RAND_303[7:0];
  _RAND_304 = {1{`RANDOM}};
  lineBuffer_297 = _RAND_304[7:0];
  _RAND_305 = {1{`RANDOM}};
  lineBuffer_298 = _RAND_305[7:0];
  _RAND_306 = {1{`RANDOM}};
  lineBuffer_299 = _RAND_306[7:0];
  _RAND_307 = {1{`RANDOM}};
  lineBuffer_300 = _RAND_307[7:0];
  _RAND_308 = {1{`RANDOM}};
  lineBuffer_301 = _RAND_308[7:0];
  _RAND_309 = {1{`RANDOM}};
  lineBuffer_302 = _RAND_309[7:0];
  _RAND_310 = {1{`RANDOM}};
  lineBuffer_303 = _RAND_310[7:0];
  _RAND_311 = {1{`RANDOM}};
  lineBuffer_304 = _RAND_311[7:0];
  _RAND_312 = {1{`RANDOM}};
  lineBuffer_305 = _RAND_312[7:0];
  _RAND_313 = {1{`RANDOM}};
  lineBuffer_306 = _RAND_313[7:0];
  _RAND_314 = {1{`RANDOM}};
  lineBuffer_307 = _RAND_314[7:0];
  _RAND_315 = {1{`RANDOM}};
  lineBuffer_308 = _RAND_315[7:0];
  _RAND_316 = {1{`RANDOM}};
  lineBuffer_309 = _RAND_316[7:0];
  _RAND_317 = {1{`RANDOM}};
  lineBuffer_310 = _RAND_317[7:0];
  _RAND_318 = {1{`RANDOM}};
  lineBuffer_311 = _RAND_318[7:0];
  _RAND_319 = {1{`RANDOM}};
  lineBuffer_312 = _RAND_319[7:0];
  _RAND_320 = {1{`RANDOM}};
  lineBuffer_313 = _RAND_320[7:0];
  _RAND_321 = {1{`RANDOM}};
  lineBuffer_314 = _RAND_321[7:0];
  _RAND_322 = {1{`RANDOM}};
  lineBuffer_315 = _RAND_322[7:0];
  _RAND_323 = {1{`RANDOM}};
  lineBuffer_316 = _RAND_323[7:0];
  _RAND_324 = {1{`RANDOM}};
  lineBuffer_317 = _RAND_324[7:0];
  _RAND_325 = {1{`RANDOM}};
  lineBuffer_318 = _RAND_325[7:0];
  _RAND_326 = {1{`RANDOM}};
  lineBuffer_319 = _RAND_326[7:0];
  _RAND_327 = {1{`RANDOM}};
  lineBuffer_320 = _RAND_327[7:0];
  _RAND_328 = {1{`RANDOM}};
  lineBuffer_321 = _RAND_328[7:0];
  _RAND_329 = {1{`RANDOM}};
  lineBuffer_322 = _RAND_329[7:0];
  _RAND_330 = {1{`RANDOM}};
  lineBuffer_323 = _RAND_330[7:0];
  _RAND_331 = {1{`RANDOM}};
  lineBuffer_324 = _RAND_331[7:0];
  _RAND_332 = {1{`RANDOM}};
  lineBuffer_325 = _RAND_332[7:0];
  _RAND_333 = {1{`RANDOM}};
  lineBuffer_326 = _RAND_333[7:0];
  _RAND_334 = {1{`RANDOM}};
  lineBuffer_327 = _RAND_334[7:0];
  _RAND_335 = {1{`RANDOM}};
  lineBuffer_328 = _RAND_335[7:0];
  _RAND_336 = {1{`RANDOM}};
  lineBuffer_329 = _RAND_336[7:0];
  _RAND_337 = {1{`RANDOM}};
  lineBuffer_330 = _RAND_337[7:0];
  _RAND_338 = {1{`RANDOM}};
  lineBuffer_331 = _RAND_338[7:0];
  _RAND_339 = {1{`RANDOM}};
  lineBuffer_332 = _RAND_339[7:0];
  _RAND_340 = {1{`RANDOM}};
  lineBuffer_333 = _RAND_340[7:0];
  _RAND_341 = {1{`RANDOM}};
  lineBuffer_334 = _RAND_341[7:0];
  _RAND_342 = {1{`RANDOM}};
  lineBuffer_335 = _RAND_342[7:0];
  _RAND_343 = {1{`RANDOM}};
  lineBuffer_336 = _RAND_343[7:0];
  _RAND_344 = {1{`RANDOM}};
  lineBuffer_337 = _RAND_344[7:0];
  _RAND_345 = {1{`RANDOM}};
  lineBuffer_338 = _RAND_345[7:0];
  _RAND_346 = {1{`RANDOM}};
  lineBuffer_339 = _RAND_346[7:0];
  _RAND_347 = {1{`RANDOM}};
  lineBuffer_340 = _RAND_347[7:0];
  _RAND_348 = {1{`RANDOM}};
  lineBuffer_341 = _RAND_348[7:0];
  _RAND_349 = {1{`RANDOM}};
  lineBuffer_342 = _RAND_349[7:0];
  _RAND_350 = {1{`RANDOM}};
  lineBuffer_343 = _RAND_350[7:0];
  _RAND_351 = {1{`RANDOM}};
  lineBuffer_344 = _RAND_351[7:0];
  _RAND_352 = {1{`RANDOM}};
  lineBuffer_345 = _RAND_352[7:0];
  _RAND_353 = {1{`RANDOM}};
  lineBuffer_346 = _RAND_353[7:0];
  _RAND_354 = {1{`RANDOM}};
  lineBuffer_347 = _RAND_354[7:0];
  _RAND_355 = {1{`RANDOM}};
  lineBuffer_348 = _RAND_355[7:0];
  _RAND_356 = {1{`RANDOM}};
  lineBuffer_349 = _RAND_356[7:0];
  _RAND_357 = {1{`RANDOM}};
  lineBuffer_350 = _RAND_357[7:0];
  _RAND_358 = {1{`RANDOM}};
  lineBuffer_351 = _RAND_358[7:0];
  _RAND_359 = {1{`RANDOM}};
  lineBuffer_352 = _RAND_359[7:0];
  _RAND_360 = {1{`RANDOM}};
  lineBuffer_353 = _RAND_360[7:0];
  _RAND_361 = {1{`RANDOM}};
  lineBuffer_354 = _RAND_361[7:0];
  _RAND_362 = {1{`RANDOM}};
  lineBuffer_355 = _RAND_362[7:0];
  _RAND_363 = {1{`RANDOM}};
  lineBuffer_356 = _RAND_363[7:0];
  _RAND_364 = {1{`RANDOM}};
  lineBuffer_357 = _RAND_364[7:0];
  _RAND_365 = {1{`RANDOM}};
  lineBuffer_358 = _RAND_365[7:0];
  _RAND_366 = {1{`RANDOM}};
  lineBuffer_359 = _RAND_366[7:0];
  _RAND_367 = {1{`RANDOM}};
  lineBuffer_360 = _RAND_367[7:0];
  _RAND_368 = {1{`RANDOM}};
  lineBuffer_361 = _RAND_368[7:0];
  _RAND_369 = {1{`RANDOM}};
  lineBuffer_362 = _RAND_369[7:0];
  _RAND_370 = {1{`RANDOM}};
  lineBuffer_363 = _RAND_370[7:0];
  _RAND_371 = {1{`RANDOM}};
  lineBuffer_364 = _RAND_371[7:0];
  _RAND_372 = {1{`RANDOM}};
  lineBuffer_365 = _RAND_372[7:0];
  _RAND_373 = {1{`RANDOM}};
  lineBuffer_366 = _RAND_373[7:0];
  _RAND_374 = {1{`RANDOM}};
  lineBuffer_367 = _RAND_374[7:0];
  _RAND_375 = {1{`RANDOM}};
  lineBuffer_368 = _RAND_375[7:0];
  _RAND_376 = {1{`RANDOM}};
  lineBuffer_369 = _RAND_376[7:0];
  _RAND_377 = {1{`RANDOM}};
  lineBuffer_370 = _RAND_377[7:0];
  _RAND_378 = {1{`RANDOM}};
  lineBuffer_371 = _RAND_378[7:0];
  _RAND_379 = {1{`RANDOM}};
  lineBuffer_372 = _RAND_379[7:0];
  _RAND_380 = {1{`RANDOM}};
  lineBuffer_373 = _RAND_380[7:0];
  _RAND_381 = {1{`RANDOM}};
  lineBuffer_374 = _RAND_381[7:0];
  _RAND_382 = {1{`RANDOM}};
  lineBuffer_375 = _RAND_382[7:0];
  _RAND_383 = {1{`RANDOM}};
  lineBuffer_376 = _RAND_383[7:0];
  _RAND_384 = {1{`RANDOM}};
  lineBuffer_377 = _RAND_384[7:0];
  _RAND_385 = {1{`RANDOM}};
  lineBuffer_378 = _RAND_385[7:0];
  _RAND_386 = {1{`RANDOM}};
  lineBuffer_379 = _RAND_386[7:0];
  _RAND_387 = {1{`RANDOM}};
  lineBuffer_380 = _RAND_387[7:0];
  _RAND_388 = {1{`RANDOM}};
  lineBuffer_381 = _RAND_388[7:0];
  _RAND_389 = {1{`RANDOM}};
  lineBuffer_382 = _RAND_389[7:0];
  _RAND_390 = {1{`RANDOM}};
  lineBuffer_383 = _RAND_390[7:0];
  _RAND_391 = {1{`RANDOM}};
  lineBuffer_384 = _RAND_391[7:0];
  _RAND_392 = {1{`RANDOM}};
  lineBuffer_385 = _RAND_392[7:0];
  _RAND_393 = {1{`RANDOM}};
  lineBuffer_386 = _RAND_393[7:0];
  _RAND_394 = {1{`RANDOM}};
  lineBuffer_387 = _RAND_394[7:0];
  _RAND_395 = {1{`RANDOM}};
  lineBuffer_388 = _RAND_395[7:0];
  _RAND_396 = {1{`RANDOM}};
  lineBuffer_389 = _RAND_396[7:0];
  _RAND_397 = {1{`RANDOM}};
  lineBuffer_390 = _RAND_397[7:0];
  _RAND_398 = {1{`RANDOM}};
  lineBuffer_391 = _RAND_398[7:0];
  _RAND_399 = {1{`RANDOM}};
  lineBuffer_392 = _RAND_399[7:0];
  _RAND_400 = {1{`RANDOM}};
  lineBuffer_393 = _RAND_400[7:0];
  _RAND_401 = {1{`RANDOM}};
  lineBuffer_394 = _RAND_401[7:0];
  _RAND_402 = {1{`RANDOM}};
  lineBuffer_395 = _RAND_402[7:0];
  _RAND_403 = {1{`RANDOM}};
  lineBuffer_396 = _RAND_403[7:0];
  _RAND_404 = {1{`RANDOM}};
  lineBuffer_397 = _RAND_404[7:0];
  _RAND_405 = {1{`RANDOM}};
  lineBuffer_398 = _RAND_405[7:0];
  _RAND_406 = {1{`RANDOM}};
  lineBuffer_399 = _RAND_406[7:0];
  _RAND_407 = {1{`RANDOM}};
  lineBuffer_400 = _RAND_407[7:0];
  _RAND_408 = {1{`RANDOM}};
  lineBuffer_401 = _RAND_408[7:0];
  _RAND_409 = {1{`RANDOM}};
  lineBuffer_402 = _RAND_409[7:0];
  _RAND_410 = {1{`RANDOM}};
  lineBuffer_403 = _RAND_410[7:0];
  _RAND_411 = {1{`RANDOM}};
  lineBuffer_404 = _RAND_411[7:0];
  _RAND_412 = {1{`RANDOM}};
  lineBuffer_405 = _RAND_412[7:0];
  _RAND_413 = {1{`RANDOM}};
  lineBuffer_406 = _RAND_413[7:0];
  _RAND_414 = {1{`RANDOM}};
  lineBuffer_407 = _RAND_414[7:0];
  _RAND_415 = {1{`RANDOM}};
  lineBuffer_408 = _RAND_415[7:0];
  _RAND_416 = {1{`RANDOM}};
  lineBuffer_409 = _RAND_416[7:0];
  _RAND_417 = {1{`RANDOM}};
  lineBuffer_410 = _RAND_417[7:0];
  _RAND_418 = {1{`RANDOM}};
  lineBuffer_411 = _RAND_418[7:0];
  _RAND_419 = {1{`RANDOM}};
  lineBuffer_412 = _RAND_419[7:0];
  _RAND_420 = {1{`RANDOM}};
  lineBuffer_413 = _RAND_420[7:0];
  _RAND_421 = {1{`RANDOM}};
  lineBuffer_414 = _RAND_421[7:0];
  _RAND_422 = {1{`RANDOM}};
  lineBuffer_415 = _RAND_422[7:0];
  _RAND_423 = {1{`RANDOM}};
  lineBuffer_416 = _RAND_423[7:0];
  _RAND_424 = {1{`RANDOM}};
  lineBuffer_417 = _RAND_424[7:0];
  _RAND_425 = {1{`RANDOM}};
  lineBuffer_418 = _RAND_425[7:0];
  _RAND_426 = {1{`RANDOM}};
  lineBuffer_419 = _RAND_426[7:0];
  _RAND_427 = {1{`RANDOM}};
  lineBuffer_420 = _RAND_427[7:0];
  _RAND_428 = {1{`RANDOM}};
  lineBuffer_421 = _RAND_428[7:0];
  _RAND_429 = {1{`RANDOM}};
  lineBuffer_422 = _RAND_429[7:0];
  _RAND_430 = {1{`RANDOM}};
  lineBuffer_423 = _RAND_430[7:0];
  _RAND_431 = {1{`RANDOM}};
  lineBuffer_424 = _RAND_431[7:0];
  _RAND_432 = {1{`RANDOM}};
  lineBuffer_425 = _RAND_432[7:0];
  _RAND_433 = {1{`RANDOM}};
  lineBuffer_426 = _RAND_433[7:0];
  _RAND_434 = {1{`RANDOM}};
  lineBuffer_427 = _RAND_434[7:0];
  _RAND_435 = {1{`RANDOM}};
  lineBuffer_428 = _RAND_435[7:0];
  _RAND_436 = {1{`RANDOM}};
  lineBuffer_429 = _RAND_436[7:0];
  _RAND_437 = {1{`RANDOM}};
  lineBuffer_430 = _RAND_437[7:0];
  _RAND_438 = {1{`RANDOM}};
  lineBuffer_431 = _RAND_438[7:0];
  _RAND_439 = {1{`RANDOM}};
  lineBuffer_432 = _RAND_439[7:0];
  _RAND_440 = {1{`RANDOM}};
  lineBuffer_433 = _RAND_440[7:0];
  _RAND_441 = {1{`RANDOM}};
  lineBuffer_434 = _RAND_441[7:0];
  _RAND_442 = {1{`RANDOM}};
  lineBuffer_435 = _RAND_442[7:0];
  _RAND_443 = {1{`RANDOM}};
  lineBuffer_436 = _RAND_443[7:0];
  _RAND_444 = {1{`RANDOM}};
  lineBuffer_437 = _RAND_444[7:0];
  _RAND_445 = {1{`RANDOM}};
  lineBuffer_438 = _RAND_445[7:0];
  _RAND_446 = {1{`RANDOM}};
  lineBuffer_439 = _RAND_446[7:0];
  _RAND_447 = {1{`RANDOM}};
  lineBuffer_440 = _RAND_447[7:0];
  _RAND_448 = {1{`RANDOM}};
  lineBuffer_441 = _RAND_448[7:0];
  _RAND_449 = {1{`RANDOM}};
  lineBuffer_442 = _RAND_449[7:0];
  _RAND_450 = {1{`RANDOM}};
  lineBuffer_443 = _RAND_450[7:0];
  _RAND_451 = {1{`RANDOM}};
  lineBuffer_444 = _RAND_451[7:0];
  _RAND_452 = {1{`RANDOM}};
  lineBuffer_445 = _RAND_452[7:0];
  _RAND_453 = {1{`RANDOM}};
  lineBuffer_446 = _RAND_453[7:0];
  _RAND_454 = {1{`RANDOM}};
  lineBuffer_447 = _RAND_454[7:0];
  _RAND_455 = {1{`RANDOM}};
  lineBuffer_448 = _RAND_455[7:0];
  _RAND_456 = {1{`RANDOM}};
  lineBuffer_449 = _RAND_456[7:0];
  _RAND_457 = {1{`RANDOM}};
  lineBuffer_450 = _RAND_457[7:0];
  _RAND_458 = {1{`RANDOM}};
  lineBuffer_451 = _RAND_458[7:0];
  _RAND_459 = {1{`RANDOM}};
  lineBuffer_452 = _RAND_459[7:0];
  _RAND_460 = {1{`RANDOM}};
  lineBuffer_453 = _RAND_460[7:0];
  _RAND_461 = {1{`RANDOM}};
  lineBuffer_454 = _RAND_461[7:0];
  _RAND_462 = {1{`RANDOM}};
  lineBuffer_455 = _RAND_462[7:0];
  _RAND_463 = {1{`RANDOM}};
  lineBuffer_456 = _RAND_463[7:0];
  _RAND_464 = {1{`RANDOM}};
  lineBuffer_457 = _RAND_464[7:0];
  _RAND_465 = {1{`RANDOM}};
  lineBuffer_458 = _RAND_465[7:0];
  _RAND_466 = {1{`RANDOM}};
  lineBuffer_459 = _RAND_466[7:0];
  _RAND_467 = {1{`RANDOM}};
  lineBuffer_460 = _RAND_467[7:0];
  _RAND_468 = {1{`RANDOM}};
  lineBuffer_461 = _RAND_468[7:0];
  _RAND_469 = {1{`RANDOM}};
  lineBuffer_462 = _RAND_469[7:0];
  _RAND_470 = {1{`RANDOM}};
  lineBuffer_463 = _RAND_470[7:0];
  _RAND_471 = {1{`RANDOM}};
  lineBuffer_464 = _RAND_471[7:0];
  _RAND_472 = {1{`RANDOM}};
  lineBuffer_465 = _RAND_472[7:0];
  _RAND_473 = {1{`RANDOM}};
  lineBuffer_466 = _RAND_473[7:0];
  _RAND_474 = {1{`RANDOM}};
  lineBuffer_467 = _RAND_474[7:0];
  _RAND_475 = {1{`RANDOM}};
  lineBuffer_468 = _RAND_475[7:0];
  _RAND_476 = {1{`RANDOM}};
  lineBuffer_469 = _RAND_476[7:0];
  _RAND_477 = {1{`RANDOM}};
  lineBuffer_470 = _RAND_477[7:0];
  _RAND_478 = {1{`RANDOM}};
  lineBuffer_471 = _RAND_478[7:0];
  _RAND_479 = {1{`RANDOM}};
  lineBuffer_472 = _RAND_479[7:0];
  _RAND_480 = {1{`RANDOM}};
  lineBuffer_473 = _RAND_480[7:0];
  _RAND_481 = {1{`RANDOM}};
  lineBuffer_474 = _RAND_481[7:0];
  _RAND_482 = {1{`RANDOM}};
  lineBuffer_475 = _RAND_482[7:0];
  _RAND_483 = {1{`RANDOM}};
  lineBuffer_476 = _RAND_483[7:0];
  _RAND_484 = {1{`RANDOM}};
  lineBuffer_477 = _RAND_484[7:0];
  _RAND_485 = {1{`RANDOM}};
  lineBuffer_478 = _RAND_485[7:0];
  _RAND_486 = {1{`RANDOM}};
  lineBuffer_479 = _RAND_486[7:0];
  _RAND_487 = {1{`RANDOM}};
  lineBuffer_480 = _RAND_487[7:0];
  _RAND_488 = {1{`RANDOM}};
  lineBuffer_481 = _RAND_488[7:0];
  _RAND_489 = {1{`RANDOM}};
  lineBuffer_482 = _RAND_489[7:0];
  _RAND_490 = {1{`RANDOM}};
  lineBuffer_483 = _RAND_490[7:0];
  _RAND_491 = {1{`RANDOM}};
  lineBuffer_484 = _RAND_491[7:0];
  _RAND_492 = {1{`RANDOM}};
  lineBuffer_485 = _RAND_492[7:0];
  _RAND_493 = {1{`RANDOM}};
  lineBuffer_486 = _RAND_493[7:0];
  _RAND_494 = {1{`RANDOM}};
  lineBuffer_487 = _RAND_494[7:0];
  _RAND_495 = {1{`RANDOM}};
  lineBuffer_488 = _RAND_495[7:0];
  _RAND_496 = {1{`RANDOM}};
  lineBuffer_489 = _RAND_496[7:0];
  _RAND_497 = {1{`RANDOM}};
  lineBuffer_490 = _RAND_497[7:0];
  _RAND_498 = {1{`RANDOM}};
  lineBuffer_491 = _RAND_498[7:0];
  _RAND_499 = {1{`RANDOM}};
  lineBuffer_492 = _RAND_499[7:0];
  _RAND_500 = {1{`RANDOM}};
  lineBuffer_493 = _RAND_500[7:0];
  _RAND_501 = {1{`RANDOM}};
  lineBuffer_494 = _RAND_501[7:0];
  _RAND_502 = {1{`RANDOM}};
  lineBuffer_495 = _RAND_502[7:0];
  _RAND_503 = {1{`RANDOM}};
  lineBuffer_496 = _RAND_503[7:0];
  _RAND_504 = {1{`RANDOM}};
  lineBuffer_497 = _RAND_504[7:0];
  _RAND_505 = {1{`RANDOM}};
  lineBuffer_498 = _RAND_505[7:0];
  _RAND_506 = {1{`RANDOM}};
  lineBuffer_499 = _RAND_506[7:0];
  _RAND_507 = {1{`RANDOM}};
  lineBuffer_500 = _RAND_507[7:0];
  _RAND_508 = {1{`RANDOM}};
  lineBuffer_501 = _RAND_508[7:0];
  _RAND_509 = {1{`RANDOM}};
  lineBuffer_502 = _RAND_509[7:0];
  _RAND_510 = {1{`RANDOM}};
  lineBuffer_503 = _RAND_510[7:0];
  _RAND_511 = {1{`RANDOM}};
  lineBuffer_504 = _RAND_511[7:0];
  _RAND_512 = {1{`RANDOM}};
  lineBuffer_505 = _RAND_512[7:0];
  _RAND_513 = {1{`RANDOM}};
  lineBuffer_506 = _RAND_513[7:0];
  _RAND_514 = {1{`RANDOM}};
  lineBuffer_507 = _RAND_514[7:0];
  _RAND_515 = {1{`RANDOM}};
  lineBuffer_508 = _RAND_515[7:0];
  _RAND_516 = {1{`RANDOM}};
  lineBuffer_509 = _RAND_516[7:0];
  _RAND_517 = {1{`RANDOM}};
  lineBuffer_510 = _RAND_517[7:0];
  _RAND_518 = {1{`RANDOM}};
  lineBuffer_511 = _RAND_518[7:0];
  _RAND_519 = {1{`RANDOM}};
  lineBuffer_512 = _RAND_519[7:0];
  _RAND_520 = {1{`RANDOM}};
  lineBuffer_513 = _RAND_520[7:0];
  _RAND_521 = {1{`RANDOM}};
  lineBuffer_514 = _RAND_521[7:0];
  _RAND_522 = {1{`RANDOM}};
  lineBuffer_515 = _RAND_522[7:0];
  _RAND_523 = {1{`RANDOM}};
  lineBuffer_516 = _RAND_523[7:0];
  _RAND_524 = {1{`RANDOM}};
  lineBuffer_517 = _RAND_524[7:0];
  _RAND_525 = {1{`RANDOM}};
  lineBuffer_518 = _RAND_525[7:0];
  _RAND_526 = {1{`RANDOM}};
  lineBuffer_519 = _RAND_526[7:0];
  _RAND_527 = {1{`RANDOM}};
  lineBuffer_520 = _RAND_527[7:0];
  _RAND_528 = {1{`RANDOM}};
  lineBuffer_521 = _RAND_528[7:0];
  _RAND_529 = {1{`RANDOM}};
  lineBuffer_522 = _RAND_529[7:0];
  _RAND_530 = {1{`RANDOM}};
  lineBuffer_523 = _RAND_530[7:0];
  _RAND_531 = {1{`RANDOM}};
  lineBuffer_524 = _RAND_531[7:0];
  _RAND_532 = {1{`RANDOM}};
  lineBuffer_525 = _RAND_532[7:0];
  _RAND_533 = {1{`RANDOM}};
  lineBuffer_526 = _RAND_533[7:0];
  _RAND_534 = {1{`RANDOM}};
  lineBuffer_527 = _RAND_534[7:0];
  _RAND_535 = {1{`RANDOM}};
  lineBuffer_528 = _RAND_535[7:0];
  _RAND_536 = {1{`RANDOM}};
  lineBuffer_529 = _RAND_536[7:0];
  _RAND_537 = {1{`RANDOM}};
  lineBuffer_530 = _RAND_537[7:0];
  _RAND_538 = {1{`RANDOM}};
  lineBuffer_531 = _RAND_538[7:0];
  _RAND_539 = {1{`RANDOM}};
  lineBuffer_532 = _RAND_539[7:0];
  _RAND_540 = {1{`RANDOM}};
  lineBuffer_533 = _RAND_540[7:0];
  _RAND_541 = {1{`RANDOM}};
  lineBuffer_534 = _RAND_541[7:0];
  _RAND_542 = {1{`RANDOM}};
  lineBuffer_535 = _RAND_542[7:0];
  _RAND_543 = {1{`RANDOM}};
  lineBuffer_536 = _RAND_543[7:0];
  _RAND_544 = {1{`RANDOM}};
  lineBuffer_537 = _RAND_544[7:0];
  _RAND_545 = {1{`RANDOM}};
  lineBuffer_538 = _RAND_545[7:0];
  _RAND_546 = {1{`RANDOM}};
  lineBuffer_539 = _RAND_546[7:0];
  _RAND_547 = {1{`RANDOM}};
  lineBuffer_540 = _RAND_547[7:0];
  _RAND_548 = {1{`RANDOM}};
  lineBuffer_541 = _RAND_548[7:0];
  _RAND_549 = {1{`RANDOM}};
  lineBuffer_542 = _RAND_549[7:0];
  _RAND_550 = {1{`RANDOM}};
  lineBuffer_543 = _RAND_550[7:0];
  _RAND_551 = {1{`RANDOM}};
  lineBuffer_544 = _RAND_551[7:0];
  _RAND_552 = {1{`RANDOM}};
  lineBuffer_545 = _RAND_552[7:0];
  _RAND_553 = {1{`RANDOM}};
  lineBuffer_546 = _RAND_553[7:0];
  _RAND_554 = {1{`RANDOM}};
  lineBuffer_547 = _RAND_554[7:0];
  _RAND_555 = {1{`RANDOM}};
  lineBuffer_548 = _RAND_555[7:0];
  _RAND_556 = {1{`RANDOM}};
  lineBuffer_549 = _RAND_556[7:0];
  _RAND_557 = {1{`RANDOM}};
  lineBuffer_550 = _RAND_557[7:0];
  _RAND_558 = {1{`RANDOM}};
  lineBuffer_551 = _RAND_558[7:0];
  _RAND_559 = {1{`RANDOM}};
  lineBuffer_552 = _RAND_559[7:0];
  _RAND_560 = {1{`RANDOM}};
  lineBuffer_553 = _RAND_560[7:0];
  _RAND_561 = {1{`RANDOM}};
  lineBuffer_554 = _RAND_561[7:0];
  _RAND_562 = {1{`RANDOM}};
  lineBuffer_555 = _RAND_562[7:0];
  _RAND_563 = {1{`RANDOM}};
  lineBuffer_556 = _RAND_563[7:0];
  _RAND_564 = {1{`RANDOM}};
  lineBuffer_557 = _RAND_564[7:0];
  _RAND_565 = {1{`RANDOM}};
  lineBuffer_558 = _RAND_565[7:0];
  _RAND_566 = {1{`RANDOM}};
  lineBuffer_559 = _RAND_566[7:0];
  _RAND_567 = {1{`RANDOM}};
  lineBuffer_560 = _RAND_567[7:0];
  _RAND_568 = {1{`RANDOM}};
  lineBuffer_561 = _RAND_568[7:0];
  _RAND_569 = {1{`RANDOM}};
  lineBuffer_562 = _RAND_569[7:0];
  _RAND_570 = {1{`RANDOM}};
  lineBuffer_563 = _RAND_570[7:0];
  _RAND_571 = {1{`RANDOM}};
  lineBuffer_564 = _RAND_571[7:0];
  _RAND_572 = {1{`RANDOM}};
  lineBuffer_565 = _RAND_572[7:0];
  _RAND_573 = {1{`RANDOM}};
  lineBuffer_566 = _RAND_573[7:0];
  _RAND_574 = {1{`RANDOM}};
  lineBuffer_567 = _RAND_574[7:0];
  _RAND_575 = {1{`RANDOM}};
  lineBuffer_568 = _RAND_575[7:0];
  _RAND_576 = {1{`RANDOM}};
  lineBuffer_569 = _RAND_576[7:0];
  _RAND_577 = {1{`RANDOM}};
  lineBuffer_570 = _RAND_577[7:0];
  _RAND_578 = {1{`RANDOM}};
  lineBuffer_571 = _RAND_578[7:0];
  _RAND_579 = {1{`RANDOM}};
  lineBuffer_572 = _RAND_579[7:0];
  _RAND_580 = {1{`RANDOM}};
  lineBuffer_573 = _RAND_580[7:0];
  _RAND_581 = {1{`RANDOM}};
  lineBuffer_574 = _RAND_581[7:0];
  _RAND_582 = {1{`RANDOM}};
  lineBuffer_575 = _RAND_582[7:0];
  _RAND_583 = {1{`RANDOM}};
  lineBuffer_576 = _RAND_583[7:0];
  _RAND_584 = {1{`RANDOM}};
  lineBuffer_577 = _RAND_584[7:0];
  _RAND_585 = {1{`RANDOM}};
  lineBuffer_578 = _RAND_585[7:0];
  _RAND_586 = {1{`RANDOM}};
  lineBuffer_579 = _RAND_586[7:0];
  _RAND_587 = {1{`RANDOM}};
  lineBuffer_580 = _RAND_587[7:0];
  _RAND_588 = {1{`RANDOM}};
  lineBuffer_581 = _RAND_588[7:0];
  _RAND_589 = {1{`RANDOM}};
  lineBuffer_582 = _RAND_589[7:0];
  _RAND_590 = {1{`RANDOM}};
  lineBuffer_583 = _RAND_590[7:0];
  _RAND_591 = {1{`RANDOM}};
  lineBuffer_584 = _RAND_591[7:0];
  _RAND_592 = {1{`RANDOM}};
  lineBuffer_585 = _RAND_592[7:0];
  _RAND_593 = {1{`RANDOM}};
  lineBuffer_586 = _RAND_593[7:0];
  _RAND_594 = {1{`RANDOM}};
  lineBuffer_587 = _RAND_594[7:0];
  _RAND_595 = {1{`RANDOM}};
  lineBuffer_588 = _RAND_595[7:0];
  _RAND_596 = {1{`RANDOM}};
  lineBuffer_589 = _RAND_596[7:0];
  _RAND_597 = {1{`RANDOM}};
  lineBuffer_590 = _RAND_597[7:0];
  _RAND_598 = {1{`RANDOM}};
  lineBuffer_591 = _RAND_598[7:0];
  _RAND_599 = {1{`RANDOM}};
  lineBuffer_592 = _RAND_599[7:0];
  _RAND_600 = {1{`RANDOM}};
  lineBuffer_593 = _RAND_600[7:0];
  _RAND_601 = {1{`RANDOM}};
  lineBuffer_594 = _RAND_601[7:0];
  _RAND_602 = {1{`RANDOM}};
  lineBuffer_595 = _RAND_602[7:0];
  _RAND_603 = {1{`RANDOM}};
  lineBuffer_596 = _RAND_603[7:0];
  _RAND_604 = {1{`RANDOM}};
  lineBuffer_597 = _RAND_604[7:0];
  _RAND_605 = {1{`RANDOM}};
  lineBuffer_598 = _RAND_605[7:0];
  _RAND_606 = {1{`RANDOM}};
  lineBuffer_599 = _RAND_606[7:0];
  _RAND_607 = {1{`RANDOM}};
  lineBuffer_600 = _RAND_607[7:0];
  _RAND_608 = {1{`RANDOM}};
  lineBuffer_601 = _RAND_608[7:0];
  _RAND_609 = {1{`RANDOM}};
  lineBuffer_602 = _RAND_609[7:0];
  _RAND_610 = {1{`RANDOM}};
  lineBuffer_603 = _RAND_610[7:0];
  _RAND_611 = {1{`RANDOM}};
  lineBuffer_604 = _RAND_611[7:0];
  _RAND_612 = {1{`RANDOM}};
  lineBuffer_605 = _RAND_612[7:0];
  _RAND_613 = {1{`RANDOM}};
  lineBuffer_606 = _RAND_613[7:0];
  _RAND_614 = {1{`RANDOM}};
  lineBuffer_607 = _RAND_614[7:0];
  _RAND_615 = {1{`RANDOM}};
  lineBuffer_608 = _RAND_615[7:0];
  _RAND_616 = {1{`RANDOM}};
  lineBuffer_609 = _RAND_616[7:0];
  _RAND_617 = {1{`RANDOM}};
  lineBuffer_610 = _RAND_617[7:0];
  _RAND_618 = {1{`RANDOM}};
  lineBuffer_611 = _RAND_618[7:0];
  _RAND_619 = {1{`RANDOM}};
  lineBuffer_612 = _RAND_619[7:0];
  _RAND_620 = {1{`RANDOM}};
  lineBuffer_613 = _RAND_620[7:0];
  _RAND_621 = {1{`RANDOM}};
  lineBuffer_614 = _RAND_621[7:0];
  _RAND_622 = {1{`RANDOM}};
  lineBuffer_615 = _RAND_622[7:0];
  _RAND_623 = {1{`RANDOM}};
  lineBuffer_616 = _RAND_623[7:0];
  _RAND_624 = {1{`RANDOM}};
  lineBuffer_617 = _RAND_624[7:0];
  _RAND_625 = {1{`RANDOM}};
  lineBuffer_618 = _RAND_625[7:0];
  _RAND_626 = {1{`RANDOM}};
  lineBuffer_619 = _RAND_626[7:0];
  _RAND_627 = {1{`RANDOM}};
  lineBuffer_620 = _RAND_627[7:0];
  _RAND_628 = {1{`RANDOM}};
  lineBuffer_621 = _RAND_628[7:0];
  _RAND_629 = {1{`RANDOM}};
  lineBuffer_622 = _RAND_629[7:0];
  _RAND_630 = {1{`RANDOM}};
  lineBuffer_623 = _RAND_630[7:0];
  _RAND_631 = {1{`RANDOM}};
  lineBuffer_624 = _RAND_631[7:0];
  _RAND_632 = {1{`RANDOM}};
  lineBuffer_625 = _RAND_632[7:0];
  _RAND_633 = {1{`RANDOM}};
  lineBuffer_626 = _RAND_633[7:0];
  _RAND_634 = {1{`RANDOM}};
  lineBuffer_627 = _RAND_634[7:0];
  _RAND_635 = {1{`RANDOM}};
  lineBuffer_628 = _RAND_635[7:0];
  _RAND_636 = {1{`RANDOM}};
  lineBuffer_629 = _RAND_636[7:0];
  _RAND_637 = {1{`RANDOM}};
  lineBuffer_630 = _RAND_637[7:0];
  _RAND_638 = {1{`RANDOM}};
  lineBuffer_631 = _RAND_638[7:0];
  _RAND_639 = {1{`RANDOM}};
  lineBuffer_632 = _RAND_639[7:0];
  _RAND_640 = {1{`RANDOM}};
  lineBuffer_633 = _RAND_640[7:0];
  _RAND_641 = {1{`RANDOM}};
  lineBuffer_634 = _RAND_641[7:0];
  _RAND_642 = {1{`RANDOM}};
  lineBuffer_635 = _RAND_642[7:0];
  _RAND_643 = {1{`RANDOM}};
  lineBuffer_636 = _RAND_643[7:0];
  _RAND_644 = {1{`RANDOM}};
  lineBuffer_637 = _RAND_644[7:0];
  _RAND_645 = {1{`RANDOM}};
  lineBuffer_638 = _RAND_645[7:0];
  _RAND_646 = {1{`RANDOM}};
  lineBuffer_639 = _RAND_646[7:0];
  _RAND_647 = {1{`RANDOM}};
  lineBuffer_640 = _RAND_647[7:0];
  _RAND_648 = {1{`RANDOM}};
  lineBuffer_641 = _RAND_648[7:0];
  _RAND_649 = {1{`RANDOM}};
  lineBuffer_642 = _RAND_649[7:0];
  _RAND_650 = {1{`RANDOM}};
  lineBuffer_643 = _RAND_650[7:0];
  _RAND_651 = {1{`RANDOM}};
  lineBuffer_644 = _RAND_651[7:0];
  _RAND_652 = {1{`RANDOM}};
  lineBuffer_645 = _RAND_652[7:0];
  _RAND_653 = {1{`RANDOM}};
  lineBuffer_646 = _RAND_653[7:0];
  _RAND_654 = {1{`RANDOM}};
  lineBuffer_647 = _RAND_654[7:0];
  _RAND_655 = {1{`RANDOM}};
  lineBuffer_648 = _RAND_655[7:0];
  _RAND_656 = {1{`RANDOM}};
  lineBuffer_649 = _RAND_656[7:0];
  _RAND_657 = {1{`RANDOM}};
  lineBuffer_650 = _RAND_657[7:0];
  _RAND_658 = {1{`RANDOM}};
  lineBuffer_651 = _RAND_658[7:0];
  _RAND_659 = {1{`RANDOM}};
  lineBuffer_652 = _RAND_659[7:0];
  _RAND_660 = {1{`RANDOM}};
  lineBuffer_653 = _RAND_660[7:0];
  _RAND_661 = {1{`RANDOM}};
  lineBuffer_654 = _RAND_661[7:0];
  _RAND_662 = {1{`RANDOM}};
  lineBuffer_655 = _RAND_662[7:0];
  _RAND_663 = {1{`RANDOM}};
  lineBuffer_656 = _RAND_663[7:0];
  _RAND_664 = {1{`RANDOM}};
  lineBuffer_657 = _RAND_664[7:0];
  _RAND_665 = {1{`RANDOM}};
  lineBuffer_658 = _RAND_665[7:0];
  _RAND_666 = {1{`RANDOM}};
  lineBuffer_659 = _RAND_666[7:0];
  _RAND_667 = {1{`RANDOM}};
  lineBuffer_660 = _RAND_667[7:0];
  _RAND_668 = {1{`RANDOM}};
  lineBuffer_661 = _RAND_668[7:0];
  _RAND_669 = {1{`RANDOM}};
  lineBuffer_662 = _RAND_669[7:0];
  _RAND_670 = {1{`RANDOM}};
  lineBuffer_663 = _RAND_670[7:0];
  _RAND_671 = {1{`RANDOM}};
  lineBuffer_664 = _RAND_671[7:0];
  _RAND_672 = {1{`RANDOM}};
  lineBuffer_665 = _RAND_672[7:0];
  _RAND_673 = {1{`RANDOM}};
  lineBuffer_666 = _RAND_673[7:0];
  _RAND_674 = {1{`RANDOM}};
  lineBuffer_667 = _RAND_674[7:0];
  _RAND_675 = {1{`RANDOM}};
  lineBuffer_668 = _RAND_675[7:0];
  _RAND_676 = {1{`RANDOM}};
  lineBuffer_669 = _RAND_676[7:0];
  _RAND_677 = {1{`RANDOM}};
  lineBuffer_670 = _RAND_677[7:0];
  _RAND_678 = {1{`RANDOM}};
  lineBuffer_671 = _RAND_678[7:0];
  _RAND_679 = {1{`RANDOM}};
  lineBuffer_672 = _RAND_679[7:0];
  _RAND_680 = {1{`RANDOM}};
  lineBuffer_673 = _RAND_680[7:0];
  _RAND_681 = {1{`RANDOM}};
  lineBuffer_674 = _RAND_681[7:0];
  _RAND_682 = {1{`RANDOM}};
  lineBuffer_675 = _RAND_682[7:0];
  _RAND_683 = {1{`RANDOM}};
  lineBuffer_676 = _RAND_683[7:0];
  _RAND_684 = {1{`RANDOM}};
  lineBuffer_677 = _RAND_684[7:0];
  _RAND_685 = {1{`RANDOM}};
  lineBuffer_678 = _RAND_685[7:0];
  _RAND_686 = {1{`RANDOM}};
  lineBuffer_679 = _RAND_686[7:0];
  _RAND_687 = {1{`RANDOM}};
  lineBuffer_680 = _RAND_687[7:0];
  _RAND_688 = {1{`RANDOM}};
  lineBuffer_681 = _RAND_688[7:0];
  _RAND_689 = {1{`RANDOM}};
  lineBuffer_682 = _RAND_689[7:0];
  _RAND_690 = {1{`RANDOM}};
  lineBuffer_683 = _RAND_690[7:0];
  _RAND_691 = {1{`RANDOM}};
  lineBuffer_684 = _RAND_691[7:0];
  _RAND_692 = {1{`RANDOM}};
  lineBuffer_685 = _RAND_692[7:0];
  _RAND_693 = {1{`RANDOM}};
  lineBuffer_686 = _RAND_693[7:0];
  _RAND_694 = {1{`RANDOM}};
  lineBuffer_687 = _RAND_694[7:0];
  _RAND_695 = {1{`RANDOM}};
  lineBuffer_688 = _RAND_695[7:0];
  _RAND_696 = {1{`RANDOM}};
  lineBuffer_689 = _RAND_696[7:0];
  _RAND_697 = {1{`RANDOM}};
  lineBuffer_690 = _RAND_697[7:0];
  _RAND_698 = {1{`RANDOM}};
  lineBuffer_691 = _RAND_698[7:0];
  _RAND_699 = {1{`RANDOM}};
  lineBuffer_692 = _RAND_699[7:0];
  _RAND_700 = {1{`RANDOM}};
  lineBuffer_693 = _RAND_700[7:0];
  _RAND_701 = {1{`RANDOM}};
  lineBuffer_694 = _RAND_701[7:0];
  _RAND_702 = {1{`RANDOM}};
  lineBuffer_695 = _RAND_702[7:0];
  _RAND_703 = {1{`RANDOM}};
  lineBuffer_696 = _RAND_703[7:0];
  _RAND_704 = {1{`RANDOM}};
  lineBuffer_697 = _RAND_704[7:0];
  _RAND_705 = {1{`RANDOM}};
  lineBuffer_698 = _RAND_705[7:0];
  _RAND_706 = {1{`RANDOM}};
  lineBuffer_699 = _RAND_706[7:0];
  _RAND_707 = {1{`RANDOM}};
  lineBuffer_700 = _RAND_707[7:0];
  _RAND_708 = {1{`RANDOM}};
  lineBuffer_701 = _RAND_708[7:0];
  _RAND_709 = {1{`RANDOM}};
  lineBuffer_702 = _RAND_709[7:0];
  _RAND_710 = {1{`RANDOM}};
  lineBuffer_703 = _RAND_710[7:0];
  _RAND_711 = {1{`RANDOM}};
  lineBuffer_704 = _RAND_711[7:0];
  _RAND_712 = {1{`RANDOM}};
  lineBuffer_705 = _RAND_712[7:0];
  _RAND_713 = {1{`RANDOM}};
  lineBuffer_706 = _RAND_713[7:0];
  _RAND_714 = {1{`RANDOM}};
  lineBuffer_707 = _RAND_714[7:0];
  _RAND_715 = {1{`RANDOM}};
  lineBuffer_708 = _RAND_715[7:0];
  _RAND_716 = {1{`RANDOM}};
  lineBuffer_709 = _RAND_716[7:0];
  _RAND_717 = {1{`RANDOM}};
  lineBuffer_710 = _RAND_717[7:0];
  _RAND_718 = {1{`RANDOM}};
  lineBuffer_711 = _RAND_718[7:0];
  _RAND_719 = {1{`RANDOM}};
  lineBuffer_712 = _RAND_719[7:0];
  _RAND_720 = {1{`RANDOM}};
  lineBuffer_713 = _RAND_720[7:0];
  _RAND_721 = {1{`RANDOM}};
  lineBuffer_714 = _RAND_721[7:0];
  _RAND_722 = {1{`RANDOM}};
  lineBuffer_715 = _RAND_722[7:0];
  _RAND_723 = {1{`RANDOM}};
  lineBuffer_716 = _RAND_723[7:0];
  _RAND_724 = {1{`RANDOM}};
  lineBuffer_717 = _RAND_724[7:0];
  _RAND_725 = {1{`RANDOM}};
  lineBuffer_718 = _RAND_725[7:0];
  _RAND_726 = {1{`RANDOM}};
  lineBuffer_719 = _RAND_726[7:0];
  _RAND_727 = {1{`RANDOM}};
  lineBuffer_720 = _RAND_727[7:0];
  _RAND_728 = {1{`RANDOM}};
  lineBuffer_721 = _RAND_728[7:0];
  _RAND_729 = {1{`RANDOM}};
  lineBuffer_722 = _RAND_729[7:0];
  _RAND_730 = {1{`RANDOM}};
  lineBuffer_723 = _RAND_730[7:0];
  _RAND_731 = {1{`RANDOM}};
  lineBuffer_724 = _RAND_731[7:0];
  _RAND_732 = {1{`RANDOM}};
  lineBuffer_725 = _RAND_732[7:0];
  _RAND_733 = {1{`RANDOM}};
  lineBuffer_726 = _RAND_733[7:0];
  _RAND_734 = {1{`RANDOM}};
  lineBuffer_727 = _RAND_734[7:0];
  _RAND_735 = {1{`RANDOM}};
  lineBuffer_728 = _RAND_735[7:0];
  _RAND_736 = {1{`RANDOM}};
  lineBuffer_729 = _RAND_736[7:0];
  _RAND_737 = {1{`RANDOM}};
  lineBuffer_730 = _RAND_737[7:0];
  _RAND_738 = {1{`RANDOM}};
  lineBuffer_731 = _RAND_738[7:0];
  _RAND_739 = {1{`RANDOM}};
  lineBuffer_732 = _RAND_739[7:0];
  _RAND_740 = {1{`RANDOM}};
  lineBuffer_733 = _RAND_740[7:0];
  _RAND_741 = {1{`RANDOM}};
  lineBuffer_734 = _RAND_741[7:0];
  _RAND_742 = {1{`RANDOM}};
  lineBuffer_735 = _RAND_742[7:0];
  _RAND_743 = {1{`RANDOM}};
  lineBuffer_736 = _RAND_743[7:0];
  _RAND_744 = {1{`RANDOM}};
  lineBuffer_737 = _RAND_744[7:0];
  _RAND_745 = {1{`RANDOM}};
  lineBuffer_738 = _RAND_745[7:0];
  _RAND_746 = {1{`RANDOM}};
  lineBuffer_739 = _RAND_746[7:0];
  _RAND_747 = {1{`RANDOM}};
  lineBuffer_740 = _RAND_747[7:0];
  _RAND_748 = {1{`RANDOM}};
  lineBuffer_741 = _RAND_748[7:0];
  _RAND_749 = {1{`RANDOM}};
  lineBuffer_742 = _RAND_749[7:0];
  _RAND_750 = {1{`RANDOM}};
  lineBuffer_743 = _RAND_750[7:0];
  _RAND_751 = {1{`RANDOM}};
  lineBuffer_744 = _RAND_751[7:0];
  _RAND_752 = {1{`RANDOM}};
  lineBuffer_745 = _RAND_752[7:0];
  _RAND_753 = {1{`RANDOM}};
  lineBuffer_746 = _RAND_753[7:0];
  _RAND_754 = {1{`RANDOM}};
  lineBuffer_747 = _RAND_754[7:0];
  _RAND_755 = {1{`RANDOM}};
  lineBuffer_748 = _RAND_755[7:0];
  _RAND_756 = {1{`RANDOM}};
  lineBuffer_749 = _RAND_756[7:0];
  _RAND_757 = {1{`RANDOM}};
  lineBuffer_750 = _RAND_757[7:0];
  _RAND_758 = {1{`RANDOM}};
  lineBuffer_751 = _RAND_758[7:0];
  _RAND_759 = {1{`RANDOM}};
  lineBuffer_752 = _RAND_759[7:0];
  _RAND_760 = {1{`RANDOM}};
  lineBuffer_753 = _RAND_760[7:0];
  _RAND_761 = {1{`RANDOM}};
  lineBuffer_754 = _RAND_761[7:0];
  _RAND_762 = {1{`RANDOM}};
  lineBuffer_755 = _RAND_762[7:0];
  _RAND_763 = {1{`RANDOM}};
  lineBuffer_756 = _RAND_763[7:0];
  _RAND_764 = {1{`RANDOM}};
  lineBuffer_757 = _RAND_764[7:0];
  _RAND_765 = {1{`RANDOM}};
  lineBuffer_758 = _RAND_765[7:0];
  _RAND_766 = {1{`RANDOM}};
  lineBuffer_759 = _RAND_766[7:0];
  _RAND_767 = {1{`RANDOM}};
  lineBuffer_760 = _RAND_767[7:0];
  _RAND_768 = {1{`RANDOM}};
  lineBuffer_761 = _RAND_768[7:0];
  _RAND_769 = {1{`RANDOM}};
  lineBuffer_762 = _RAND_769[7:0];
  _RAND_770 = {1{`RANDOM}};
  lineBuffer_763 = _RAND_770[7:0];
  _RAND_771 = {1{`RANDOM}};
  lineBuffer_764 = _RAND_771[7:0];
  _RAND_772 = {1{`RANDOM}};
  lineBuffer_765 = _RAND_772[7:0];
  _RAND_773 = {1{`RANDOM}};
  lineBuffer_766 = _RAND_773[7:0];
  _RAND_774 = {1{`RANDOM}};
  lineBuffer_767 = _RAND_774[7:0];
  _RAND_775 = {1{`RANDOM}};
  lineBuffer_768 = _RAND_775[7:0];
  _RAND_776 = {1{`RANDOM}};
  lineBuffer_769 = _RAND_776[7:0];
  _RAND_777 = {1{`RANDOM}};
  lineBuffer_770 = _RAND_777[7:0];
  _RAND_778 = {1{`RANDOM}};
  lineBuffer_771 = _RAND_778[7:0];
  _RAND_779 = {1{`RANDOM}};
  lineBuffer_772 = _RAND_779[7:0];
  _RAND_780 = {1{`RANDOM}};
  lineBuffer_773 = _RAND_780[7:0];
  _RAND_781 = {1{`RANDOM}};
  lineBuffer_774 = _RAND_781[7:0];
  _RAND_782 = {1{`RANDOM}};
  lineBuffer_775 = _RAND_782[7:0];
  _RAND_783 = {1{`RANDOM}};
  lineBuffer_776 = _RAND_783[7:0];
  _RAND_784 = {1{`RANDOM}};
  lineBuffer_777 = _RAND_784[7:0];
  _RAND_785 = {1{`RANDOM}};
  lineBuffer_778 = _RAND_785[7:0];
  _RAND_786 = {1{`RANDOM}};
  lineBuffer_779 = _RAND_786[7:0];
  _RAND_787 = {1{`RANDOM}};
  lineBuffer_780 = _RAND_787[7:0];
  _RAND_788 = {1{`RANDOM}};
  lineBuffer_781 = _RAND_788[7:0];
  _RAND_789 = {1{`RANDOM}};
  lineBuffer_782 = _RAND_789[7:0];
  _RAND_790 = {1{`RANDOM}};
  lineBuffer_783 = _RAND_790[7:0];
  _RAND_791 = {1{`RANDOM}};
  lineBuffer_784 = _RAND_791[7:0];
  _RAND_792 = {1{`RANDOM}};
  lineBuffer_785 = _RAND_792[7:0];
  _RAND_793 = {1{`RANDOM}};
  lineBuffer_786 = _RAND_793[7:0];
  _RAND_794 = {1{`RANDOM}};
  lineBuffer_787 = _RAND_794[7:0];
  _RAND_795 = {1{`RANDOM}};
  lineBuffer_788 = _RAND_795[7:0];
  _RAND_796 = {1{`RANDOM}};
  lineBuffer_789 = _RAND_796[7:0];
  _RAND_797 = {1{`RANDOM}};
  lineBuffer_790 = _RAND_797[7:0];
  _RAND_798 = {1{`RANDOM}};
  lineBuffer_791 = _RAND_798[7:0];
  _RAND_799 = {1{`RANDOM}};
  lineBuffer_792 = _RAND_799[7:0];
  _RAND_800 = {1{`RANDOM}};
  lineBuffer_793 = _RAND_800[7:0];
  _RAND_801 = {1{`RANDOM}};
  lineBuffer_794 = _RAND_801[7:0];
  _RAND_802 = {1{`RANDOM}};
  lineBuffer_795 = _RAND_802[7:0];
  _RAND_803 = {1{`RANDOM}};
  lineBuffer_796 = _RAND_803[7:0];
  _RAND_804 = {1{`RANDOM}};
  lineBuffer_797 = _RAND_804[7:0];
  _RAND_805 = {1{`RANDOM}};
  lineBuffer_798 = _RAND_805[7:0];
  _RAND_806 = {1{`RANDOM}};
  lineBuffer_799 = _RAND_806[7:0];
  _RAND_807 = {1{`RANDOM}};
  lineBuffer_800 = _RAND_807[7:0];
  _RAND_808 = {1{`RANDOM}};
  lineBuffer_801 = _RAND_808[7:0];
  _RAND_809 = {1{`RANDOM}};
  lineBuffer_802 = _RAND_809[7:0];
  _RAND_810 = {1{`RANDOM}};
  lineBuffer_803 = _RAND_810[7:0];
  _RAND_811 = {1{`RANDOM}};
  lineBuffer_804 = _RAND_811[7:0];
  _RAND_812 = {1{`RANDOM}};
  lineBuffer_805 = _RAND_812[7:0];
  _RAND_813 = {1{`RANDOM}};
  lineBuffer_806 = _RAND_813[7:0];
  _RAND_814 = {1{`RANDOM}};
  lineBuffer_807 = _RAND_814[7:0];
  _RAND_815 = {1{`RANDOM}};
  lineBuffer_808 = _RAND_815[7:0];
  _RAND_816 = {1{`RANDOM}};
  lineBuffer_809 = _RAND_816[7:0];
  _RAND_817 = {1{`RANDOM}};
  lineBuffer_810 = _RAND_817[7:0];
  _RAND_818 = {1{`RANDOM}};
  lineBuffer_811 = _RAND_818[7:0];
  _RAND_819 = {1{`RANDOM}};
  lineBuffer_812 = _RAND_819[7:0];
  _RAND_820 = {1{`RANDOM}};
  lineBuffer_813 = _RAND_820[7:0];
  _RAND_821 = {1{`RANDOM}};
  lineBuffer_814 = _RAND_821[7:0];
  _RAND_822 = {1{`RANDOM}};
  lineBuffer_815 = _RAND_822[7:0];
  _RAND_823 = {1{`RANDOM}};
  lineBuffer_816 = _RAND_823[7:0];
  _RAND_824 = {1{`RANDOM}};
  lineBuffer_817 = _RAND_824[7:0];
  _RAND_825 = {1{`RANDOM}};
  lineBuffer_818 = _RAND_825[7:0];
  _RAND_826 = {1{`RANDOM}};
  lineBuffer_819 = _RAND_826[7:0];
  _RAND_827 = {1{`RANDOM}};
  lineBuffer_820 = _RAND_827[7:0];
  _RAND_828 = {1{`RANDOM}};
  lineBuffer_821 = _RAND_828[7:0];
  _RAND_829 = {1{`RANDOM}};
  lineBuffer_822 = _RAND_829[7:0];
  _RAND_830 = {1{`RANDOM}};
  lineBuffer_823 = _RAND_830[7:0];
  _RAND_831 = {1{`RANDOM}};
  lineBuffer_824 = _RAND_831[7:0];
  _RAND_832 = {1{`RANDOM}};
  lineBuffer_825 = _RAND_832[7:0];
  _RAND_833 = {1{`RANDOM}};
  lineBuffer_826 = _RAND_833[7:0];
  _RAND_834 = {1{`RANDOM}};
  lineBuffer_827 = _RAND_834[7:0];
  _RAND_835 = {1{`RANDOM}};
  lineBuffer_828 = _RAND_835[7:0];
  _RAND_836 = {1{`RANDOM}};
  lineBuffer_829 = _RAND_836[7:0];
  _RAND_837 = {1{`RANDOM}};
  lineBuffer_830 = _RAND_837[7:0];
  _RAND_838 = {1{`RANDOM}};
  lineBuffer_831 = _RAND_838[7:0];
  _RAND_839 = {1{`RANDOM}};
  lineBuffer_832 = _RAND_839[7:0];
  _RAND_840 = {1{`RANDOM}};
  lineBuffer_833 = _RAND_840[7:0];
  _RAND_841 = {1{`RANDOM}};
  lineBuffer_834 = _RAND_841[7:0];
  _RAND_842 = {1{`RANDOM}};
  lineBuffer_835 = _RAND_842[7:0];
  _RAND_843 = {1{`RANDOM}};
  lineBuffer_836 = _RAND_843[7:0];
  _RAND_844 = {1{`RANDOM}};
  lineBuffer_837 = _RAND_844[7:0];
  _RAND_845 = {1{`RANDOM}};
  lineBuffer_838 = _RAND_845[7:0];
  _RAND_846 = {1{`RANDOM}};
  lineBuffer_839 = _RAND_846[7:0];
  _RAND_847 = {1{`RANDOM}};
  lineBuffer_840 = _RAND_847[7:0];
  _RAND_848 = {1{`RANDOM}};
  lineBuffer_841 = _RAND_848[7:0];
  _RAND_849 = {1{`RANDOM}};
  lineBuffer_842 = _RAND_849[7:0];
  _RAND_850 = {1{`RANDOM}};
  lineBuffer_843 = _RAND_850[7:0];
  _RAND_851 = {1{`RANDOM}};
  lineBuffer_844 = _RAND_851[7:0];
  _RAND_852 = {1{`RANDOM}};
  lineBuffer_845 = _RAND_852[7:0];
  _RAND_853 = {1{`RANDOM}};
  lineBuffer_846 = _RAND_853[7:0];
  _RAND_854 = {1{`RANDOM}};
  lineBuffer_847 = _RAND_854[7:0];
  _RAND_855 = {1{`RANDOM}};
  lineBuffer_848 = _RAND_855[7:0];
  _RAND_856 = {1{`RANDOM}};
  lineBuffer_849 = _RAND_856[7:0];
  _RAND_857 = {1{`RANDOM}};
  lineBuffer_850 = _RAND_857[7:0];
  _RAND_858 = {1{`RANDOM}};
  lineBuffer_851 = _RAND_858[7:0];
  _RAND_859 = {1{`RANDOM}};
  lineBuffer_852 = _RAND_859[7:0];
  _RAND_860 = {1{`RANDOM}};
  lineBuffer_853 = _RAND_860[7:0];
  _RAND_861 = {1{`RANDOM}};
  lineBuffer_854 = _RAND_861[7:0];
  _RAND_862 = {1{`RANDOM}};
  lineBuffer_855 = _RAND_862[7:0];
  _RAND_863 = {1{`RANDOM}};
  lineBuffer_856 = _RAND_863[7:0];
  _RAND_864 = {1{`RANDOM}};
  lineBuffer_857 = _RAND_864[7:0];
  _RAND_865 = {1{`RANDOM}};
  lineBuffer_858 = _RAND_865[7:0];
  _RAND_866 = {1{`RANDOM}};
  lineBuffer_859 = _RAND_866[7:0];
  _RAND_867 = {1{`RANDOM}};
  lineBuffer_860 = _RAND_867[7:0];
  _RAND_868 = {1{`RANDOM}};
  lineBuffer_861 = _RAND_868[7:0];
  _RAND_869 = {1{`RANDOM}};
  lineBuffer_862 = _RAND_869[7:0];
  _RAND_870 = {1{`RANDOM}};
  lineBuffer_863 = _RAND_870[7:0];
  _RAND_871 = {1{`RANDOM}};
  lineBuffer_864 = _RAND_871[7:0];
  _RAND_872 = {1{`RANDOM}};
  lineBuffer_865 = _RAND_872[7:0];
  _RAND_873 = {1{`RANDOM}};
  lineBuffer_866 = _RAND_873[7:0];
  _RAND_874 = {1{`RANDOM}};
  lineBuffer_867 = _RAND_874[7:0];
  _RAND_875 = {1{`RANDOM}};
  lineBuffer_868 = _RAND_875[7:0];
  _RAND_876 = {1{`RANDOM}};
  lineBuffer_869 = _RAND_876[7:0];
  _RAND_877 = {1{`RANDOM}};
  lineBuffer_870 = _RAND_877[7:0];
  _RAND_878 = {1{`RANDOM}};
  lineBuffer_871 = _RAND_878[7:0];
  _RAND_879 = {1{`RANDOM}};
  lineBuffer_872 = _RAND_879[7:0];
  _RAND_880 = {1{`RANDOM}};
  lineBuffer_873 = _RAND_880[7:0];
  _RAND_881 = {1{`RANDOM}};
  lineBuffer_874 = _RAND_881[7:0];
  _RAND_882 = {1{`RANDOM}};
  lineBuffer_875 = _RAND_882[7:0];
  _RAND_883 = {1{`RANDOM}};
  lineBuffer_876 = _RAND_883[7:0];
  _RAND_884 = {1{`RANDOM}};
  lineBuffer_877 = _RAND_884[7:0];
  _RAND_885 = {1{`RANDOM}};
  lineBuffer_878 = _RAND_885[7:0];
  _RAND_886 = {1{`RANDOM}};
  lineBuffer_879 = _RAND_886[7:0];
  _RAND_887 = {1{`RANDOM}};
  lineBuffer_880 = _RAND_887[7:0];
  _RAND_888 = {1{`RANDOM}};
  lineBuffer_881 = _RAND_888[7:0];
  _RAND_889 = {1{`RANDOM}};
  lineBuffer_882 = _RAND_889[7:0];
  _RAND_890 = {1{`RANDOM}};
  lineBuffer_883 = _RAND_890[7:0];
  _RAND_891 = {1{`RANDOM}};
  lineBuffer_884 = _RAND_891[7:0];
  _RAND_892 = {1{`RANDOM}};
  lineBuffer_885 = _RAND_892[7:0];
  _RAND_893 = {1{`RANDOM}};
  lineBuffer_886 = _RAND_893[7:0];
  _RAND_894 = {1{`RANDOM}};
  lineBuffer_887 = _RAND_894[7:0];
  _RAND_895 = {1{`RANDOM}};
  lineBuffer_888 = _RAND_895[7:0];
  _RAND_896 = {1{`RANDOM}};
  lineBuffer_889 = _RAND_896[7:0];
  _RAND_897 = {1{`RANDOM}};
  lineBuffer_890 = _RAND_897[7:0];
  _RAND_898 = {1{`RANDOM}};
  lineBuffer_891 = _RAND_898[7:0];
  _RAND_899 = {1{`RANDOM}};
  lineBuffer_892 = _RAND_899[7:0];
  _RAND_900 = {1{`RANDOM}};
  lineBuffer_893 = _RAND_900[7:0];
  _RAND_901 = {1{`RANDOM}};
  lineBuffer_894 = _RAND_901[7:0];
  _RAND_902 = {1{`RANDOM}};
  lineBuffer_895 = _RAND_902[7:0];
  _RAND_903 = {1{`RANDOM}};
  lineBuffer_896 = _RAND_903[7:0];
  _RAND_904 = {1{`RANDOM}};
  lineBuffer_897 = _RAND_904[7:0];
  _RAND_905 = {1{`RANDOM}};
  lineBuffer_898 = _RAND_905[7:0];
  _RAND_906 = {1{`RANDOM}};
  lineBuffer_899 = _RAND_906[7:0];
  _RAND_907 = {1{`RANDOM}};
  lineBuffer_900 = _RAND_907[7:0];
  _RAND_908 = {1{`RANDOM}};
  lineBuffer_901 = _RAND_908[7:0];
  _RAND_909 = {1{`RANDOM}};
  lineBuffer_902 = _RAND_909[7:0];
  _RAND_910 = {1{`RANDOM}};
  lineBuffer_903 = _RAND_910[7:0];
  _RAND_911 = {1{`RANDOM}};
  lineBuffer_904 = _RAND_911[7:0];
  _RAND_912 = {1{`RANDOM}};
  lineBuffer_905 = _RAND_912[7:0];
  _RAND_913 = {1{`RANDOM}};
  lineBuffer_906 = _RAND_913[7:0];
  _RAND_914 = {1{`RANDOM}};
  lineBuffer_907 = _RAND_914[7:0];
  _RAND_915 = {1{`RANDOM}};
  lineBuffer_908 = _RAND_915[7:0];
  _RAND_916 = {1{`RANDOM}};
  lineBuffer_909 = _RAND_916[7:0];
  _RAND_917 = {1{`RANDOM}};
  lineBuffer_910 = _RAND_917[7:0];
  _RAND_918 = {1{`RANDOM}};
  lineBuffer_911 = _RAND_918[7:0];
  _RAND_919 = {1{`RANDOM}};
  lineBuffer_912 = _RAND_919[7:0];
  _RAND_920 = {1{`RANDOM}};
  lineBuffer_913 = _RAND_920[7:0];
  _RAND_921 = {1{`RANDOM}};
  lineBuffer_914 = _RAND_921[7:0];
  _RAND_922 = {1{`RANDOM}};
  lineBuffer_915 = _RAND_922[7:0];
  _RAND_923 = {1{`RANDOM}};
  lineBuffer_916 = _RAND_923[7:0];
  _RAND_924 = {1{`RANDOM}};
  lineBuffer_917 = _RAND_924[7:0];
  _RAND_925 = {1{`RANDOM}};
  lineBuffer_918 = _RAND_925[7:0];
  _RAND_926 = {1{`RANDOM}};
  lineBuffer_919 = _RAND_926[7:0];
  _RAND_927 = {1{`RANDOM}};
  lineBuffer_920 = _RAND_927[7:0];
  _RAND_928 = {1{`RANDOM}};
  lineBuffer_921 = _RAND_928[7:0];
  _RAND_929 = {1{`RANDOM}};
  lineBuffer_922 = _RAND_929[7:0];
  _RAND_930 = {1{`RANDOM}};
  lineBuffer_923 = _RAND_930[7:0];
  _RAND_931 = {1{`RANDOM}};
  lineBuffer_924 = _RAND_931[7:0];
  _RAND_932 = {1{`RANDOM}};
  lineBuffer_925 = _RAND_932[7:0];
  _RAND_933 = {1{`RANDOM}};
  lineBuffer_926 = _RAND_933[7:0];
  _RAND_934 = {1{`RANDOM}};
  lineBuffer_927 = _RAND_934[7:0];
  _RAND_935 = {1{`RANDOM}};
  lineBuffer_928 = _RAND_935[7:0];
  _RAND_936 = {1{`RANDOM}};
  lineBuffer_929 = _RAND_936[7:0];
  _RAND_937 = {1{`RANDOM}};
  lineBuffer_930 = _RAND_937[7:0];
  _RAND_938 = {1{`RANDOM}};
  lineBuffer_931 = _RAND_938[7:0];
  _RAND_939 = {1{`RANDOM}};
  lineBuffer_932 = _RAND_939[7:0];
  _RAND_940 = {1{`RANDOM}};
  lineBuffer_933 = _RAND_940[7:0];
  _RAND_941 = {1{`RANDOM}};
  lineBuffer_934 = _RAND_941[7:0];
  _RAND_942 = {1{`RANDOM}};
  lineBuffer_935 = _RAND_942[7:0];
  _RAND_943 = {1{`RANDOM}};
  lineBuffer_936 = _RAND_943[7:0];
  _RAND_944 = {1{`RANDOM}};
  lineBuffer_937 = _RAND_944[7:0];
  _RAND_945 = {1{`RANDOM}};
  lineBuffer_938 = _RAND_945[7:0];
  _RAND_946 = {1{`RANDOM}};
  lineBuffer_939 = _RAND_946[7:0];
  _RAND_947 = {1{`RANDOM}};
  lineBuffer_940 = _RAND_947[7:0];
  _RAND_948 = {1{`RANDOM}};
  lineBuffer_941 = _RAND_948[7:0];
  _RAND_949 = {1{`RANDOM}};
  lineBuffer_942 = _RAND_949[7:0];
  _RAND_950 = {1{`RANDOM}};
  lineBuffer_943 = _RAND_950[7:0];
  _RAND_951 = {1{`RANDOM}};
  lineBuffer_944 = _RAND_951[7:0];
  _RAND_952 = {1{`RANDOM}};
  lineBuffer_945 = _RAND_952[7:0];
  _RAND_953 = {1{`RANDOM}};
  lineBuffer_946 = _RAND_953[7:0];
  _RAND_954 = {1{`RANDOM}};
  lineBuffer_947 = _RAND_954[7:0];
  _RAND_955 = {1{`RANDOM}};
  lineBuffer_948 = _RAND_955[7:0];
  _RAND_956 = {1{`RANDOM}};
  lineBuffer_949 = _RAND_956[7:0];
  _RAND_957 = {1{`RANDOM}};
  lineBuffer_950 = _RAND_957[7:0];
  _RAND_958 = {1{`RANDOM}};
  lineBuffer_951 = _RAND_958[7:0];
  _RAND_959 = {1{`RANDOM}};
  lineBuffer_952 = _RAND_959[7:0];
  _RAND_960 = {1{`RANDOM}};
  lineBuffer_953 = _RAND_960[7:0];
  _RAND_961 = {1{`RANDOM}};
  lineBuffer_954 = _RAND_961[7:0];
  _RAND_962 = {1{`RANDOM}};
  lineBuffer_955 = _RAND_962[7:0];
  _RAND_963 = {1{`RANDOM}};
  lineBuffer_956 = _RAND_963[7:0];
  _RAND_964 = {1{`RANDOM}};
  lineBuffer_957 = _RAND_964[7:0];
  _RAND_965 = {1{`RANDOM}};
  lineBuffer_958 = _RAND_965[7:0];
  _RAND_966 = {1{`RANDOM}};
  lineBuffer_959 = _RAND_966[7:0];
  _RAND_967 = {1{`RANDOM}};
  lineBuffer_960 = _RAND_967[7:0];
  _RAND_968 = {1{`RANDOM}};
  lineBuffer_961 = _RAND_968[7:0];
  _RAND_969 = {1{`RANDOM}};
  lineBuffer_962 = _RAND_969[7:0];
  _RAND_970 = {1{`RANDOM}};
  lineBuffer_963 = _RAND_970[7:0];
  _RAND_971 = {1{`RANDOM}};
  lineBuffer_964 = _RAND_971[7:0];
  _RAND_972 = {1{`RANDOM}};
  lineBuffer_965 = _RAND_972[7:0];
  _RAND_973 = {1{`RANDOM}};
  lineBuffer_966 = _RAND_973[7:0];
  _RAND_974 = {1{`RANDOM}};
  lineBuffer_967 = _RAND_974[7:0];
  _RAND_975 = {1{`RANDOM}};
  lineBuffer_968 = _RAND_975[7:0];
  _RAND_976 = {1{`RANDOM}};
  lineBuffer_969 = _RAND_976[7:0];
  _RAND_977 = {1{`RANDOM}};
  lineBuffer_970 = _RAND_977[7:0];
  _RAND_978 = {1{`RANDOM}};
  lineBuffer_971 = _RAND_978[7:0];
  _RAND_979 = {1{`RANDOM}};
  lineBuffer_972 = _RAND_979[7:0];
  _RAND_980 = {1{`RANDOM}};
  lineBuffer_973 = _RAND_980[7:0];
  _RAND_981 = {1{`RANDOM}};
  lineBuffer_974 = _RAND_981[7:0];
  _RAND_982 = {1{`RANDOM}};
  lineBuffer_975 = _RAND_982[7:0];
  _RAND_983 = {1{`RANDOM}};
  lineBuffer_976 = _RAND_983[7:0];
  _RAND_984 = {1{`RANDOM}};
  lineBuffer_977 = _RAND_984[7:0];
  _RAND_985 = {1{`RANDOM}};
  lineBuffer_978 = _RAND_985[7:0];
  _RAND_986 = {1{`RANDOM}};
  lineBuffer_979 = _RAND_986[7:0];
  _RAND_987 = {1{`RANDOM}};
  lineBuffer_980 = _RAND_987[7:0];
  _RAND_988 = {1{`RANDOM}};
  lineBuffer_981 = _RAND_988[7:0];
  _RAND_989 = {1{`RANDOM}};
  lineBuffer_982 = _RAND_989[7:0];
  _RAND_990 = {1{`RANDOM}};
  lineBuffer_983 = _RAND_990[7:0];
  _RAND_991 = {1{`RANDOM}};
  lineBuffer_984 = _RAND_991[7:0];
  _RAND_992 = {1{`RANDOM}};
  lineBuffer_985 = _RAND_992[7:0];
  _RAND_993 = {1{`RANDOM}};
  lineBuffer_986 = _RAND_993[7:0];
  _RAND_994 = {1{`RANDOM}};
  lineBuffer_987 = _RAND_994[7:0];
  _RAND_995 = {1{`RANDOM}};
  lineBuffer_988 = _RAND_995[7:0];
  _RAND_996 = {1{`RANDOM}};
  lineBuffer_989 = _RAND_996[7:0];
  _RAND_997 = {1{`RANDOM}};
  lineBuffer_990 = _RAND_997[7:0];
  _RAND_998 = {1{`RANDOM}};
  lineBuffer_991 = _RAND_998[7:0];
  _RAND_999 = {1{`RANDOM}};
  lineBuffer_992 = _RAND_999[7:0];
  _RAND_1000 = {1{`RANDOM}};
  lineBuffer_993 = _RAND_1000[7:0];
  _RAND_1001 = {1{`RANDOM}};
  lineBuffer_994 = _RAND_1001[7:0];
  _RAND_1002 = {1{`RANDOM}};
  lineBuffer_995 = _RAND_1002[7:0];
  _RAND_1003 = {1{`RANDOM}};
  lineBuffer_996 = _RAND_1003[7:0];
  _RAND_1004 = {1{`RANDOM}};
  lineBuffer_997 = _RAND_1004[7:0];
  _RAND_1005 = {1{`RANDOM}};
  lineBuffer_998 = _RAND_1005[7:0];
  _RAND_1006 = {1{`RANDOM}};
  lineBuffer_999 = _RAND_1006[7:0];
  _RAND_1007 = {1{`RANDOM}};
  lineBuffer_1000 = _RAND_1007[7:0];
  _RAND_1008 = {1{`RANDOM}};
  lineBuffer_1001 = _RAND_1008[7:0];
  _RAND_1009 = {1{`RANDOM}};
  lineBuffer_1002 = _RAND_1009[7:0];
  _RAND_1010 = {1{`RANDOM}};
  lineBuffer_1003 = _RAND_1010[7:0];
  _RAND_1011 = {1{`RANDOM}};
  lineBuffer_1004 = _RAND_1011[7:0];
  _RAND_1012 = {1{`RANDOM}};
  lineBuffer_1005 = _RAND_1012[7:0];
  _RAND_1013 = {1{`RANDOM}};
  lineBuffer_1006 = _RAND_1013[7:0];
  _RAND_1014 = {1{`RANDOM}};
  lineBuffer_1007 = _RAND_1014[7:0];
  _RAND_1015 = {1{`RANDOM}};
  lineBuffer_1008 = _RAND_1015[7:0];
  _RAND_1016 = {1{`RANDOM}};
  lineBuffer_1009 = _RAND_1016[7:0];
  _RAND_1017 = {1{`RANDOM}};
  lineBuffer_1010 = _RAND_1017[7:0];
  _RAND_1018 = {1{`RANDOM}};
  lineBuffer_1011 = _RAND_1018[7:0];
  _RAND_1019 = {1{`RANDOM}};
  lineBuffer_1012 = _RAND_1019[7:0];
  _RAND_1020 = {1{`RANDOM}};
  lineBuffer_1013 = _RAND_1020[7:0];
  _RAND_1021 = {1{`RANDOM}};
  lineBuffer_1014 = _RAND_1021[7:0];
  _RAND_1022 = {1{`RANDOM}};
  lineBuffer_1015 = _RAND_1022[7:0];
  _RAND_1023 = {1{`RANDOM}};
  lineBuffer_1016 = _RAND_1023[7:0];
  _RAND_1024 = {1{`RANDOM}};
  lineBuffer_1017 = _RAND_1024[7:0];
  _RAND_1025 = {1{`RANDOM}};
  lineBuffer_1018 = _RAND_1025[7:0];
  _RAND_1026 = {1{`RANDOM}};
  lineBuffer_1019 = _RAND_1026[7:0];
  _RAND_1027 = {1{`RANDOM}};
  lineBuffer_1020 = _RAND_1027[7:0];
  _RAND_1028 = {1{`RANDOM}};
  lineBuffer_1021 = _RAND_1028[7:0];
  _RAND_1029 = {1{`RANDOM}};
  lineBuffer_1022 = _RAND_1029[7:0];
  _RAND_1030 = {1{`RANDOM}};
  lineBuffer_1023 = _RAND_1030[7:0];
  _RAND_1031 = {1{`RANDOM}};
  lineBuffer_1024 = _RAND_1031[7:0];
  _RAND_1032 = {1{`RANDOM}};
  lineBuffer_1025 = _RAND_1032[7:0];
  _RAND_1033 = {1{`RANDOM}};
  lineBuffer_1026 = _RAND_1033[7:0];
  _RAND_1034 = {1{`RANDOM}};
  lineBuffer_1027 = _RAND_1034[7:0];
  _RAND_1035 = {1{`RANDOM}};
  lineBuffer_1028 = _RAND_1035[7:0];
  _RAND_1036 = {1{`RANDOM}};
  lineBuffer_1029 = _RAND_1036[7:0];
  _RAND_1037 = {1{`RANDOM}};
  lineBuffer_1030 = _RAND_1037[7:0];
  _RAND_1038 = {1{`RANDOM}};
  lineBuffer_1031 = _RAND_1038[7:0];
  _RAND_1039 = {1{`RANDOM}};
  lineBuffer_1032 = _RAND_1039[7:0];
  _RAND_1040 = {1{`RANDOM}};
  lineBuffer_1033 = _RAND_1040[7:0];
  _RAND_1041 = {1{`RANDOM}};
  lineBuffer_1034 = _RAND_1041[7:0];
  _RAND_1042 = {1{`RANDOM}};
  lineBuffer_1035 = _RAND_1042[7:0];
  _RAND_1043 = {1{`RANDOM}};
  lineBuffer_1036 = _RAND_1043[7:0];
  _RAND_1044 = {1{`RANDOM}};
  lineBuffer_1037 = _RAND_1044[7:0];
  _RAND_1045 = {1{`RANDOM}};
  lineBuffer_1038 = _RAND_1045[7:0];
  _RAND_1046 = {1{`RANDOM}};
  lineBuffer_1039 = _RAND_1046[7:0];
  _RAND_1047 = {1{`RANDOM}};
  lineBuffer_1040 = _RAND_1047[7:0];
  _RAND_1048 = {1{`RANDOM}};
  lineBuffer_1041 = _RAND_1048[7:0];
  _RAND_1049 = {1{`RANDOM}};
  lineBuffer_1042 = _RAND_1049[7:0];
  _RAND_1050 = {1{`RANDOM}};
  lineBuffer_1043 = _RAND_1050[7:0];
  _RAND_1051 = {1{`RANDOM}};
  lineBuffer_1044 = _RAND_1051[7:0];
  _RAND_1052 = {1{`RANDOM}};
  lineBuffer_1045 = _RAND_1052[7:0];
  _RAND_1053 = {1{`RANDOM}};
  lineBuffer_1046 = _RAND_1053[7:0];
  _RAND_1054 = {1{`RANDOM}};
  lineBuffer_1047 = _RAND_1054[7:0];
  _RAND_1055 = {1{`RANDOM}};
  lineBuffer_1048 = _RAND_1055[7:0];
  _RAND_1056 = {1{`RANDOM}};
  lineBuffer_1049 = _RAND_1056[7:0];
  _RAND_1057 = {1{`RANDOM}};
  lineBuffer_1050 = _RAND_1057[7:0];
  _RAND_1058 = {1{`RANDOM}};
  lineBuffer_1051 = _RAND_1058[7:0];
  _RAND_1059 = {1{`RANDOM}};
  lineBuffer_1052 = _RAND_1059[7:0];
  _RAND_1060 = {1{`RANDOM}};
  lineBuffer_1053 = _RAND_1060[7:0];
  _RAND_1061 = {1{`RANDOM}};
  lineBuffer_1054 = _RAND_1061[7:0];
  _RAND_1062 = {1{`RANDOM}};
  lineBuffer_1055 = _RAND_1062[7:0];
  _RAND_1063 = {1{`RANDOM}};
  lineBuffer_1056 = _RAND_1063[7:0];
  _RAND_1064 = {1{`RANDOM}};
  lineBuffer_1057 = _RAND_1064[7:0];
  _RAND_1065 = {1{`RANDOM}};
  lineBuffer_1058 = _RAND_1065[7:0];
  _RAND_1066 = {1{`RANDOM}};
  lineBuffer_1059 = _RAND_1066[7:0];
  _RAND_1067 = {1{`RANDOM}};
  lineBuffer_1060 = _RAND_1067[7:0];
  _RAND_1068 = {1{`RANDOM}};
  lineBuffer_1061 = _RAND_1068[7:0];
  _RAND_1069 = {1{`RANDOM}};
  lineBuffer_1062 = _RAND_1069[7:0];
  _RAND_1070 = {1{`RANDOM}};
  lineBuffer_1063 = _RAND_1070[7:0];
  _RAND_1071 = {1{`RANDOM}};
  lineBuffer_1064 = _RAND_1071[7:0];
  _RAND_1072 = {1{`RANDOM}};
  lineBuffer_1065 = _RAND_1072[7:0];
  _RAND_1073 = {1{`RANDOM}};
  lineBuffer_1066 = _RAND_1073[7:0];
  _RAND_1074 = {1{`RANDOM}};
  lineBuffer_1067 = _RAND_1074[7:0];
  _RAND_1075 = {1{`RANDOM}};
  lineBuffer_1068 = _RAND_1075[7:0];
  _RAND_1076 = {1{`RANDOM}};
  lineBuffer_1069 = _RAND_1076[7:0];
  _RAND_1077 = {1{`RANDOM}};
  lineBuffer_1070 = _RAND_1077[7:0];
  _RAND_1078 = {1{`RANDOM}};
  lineBuffer_1071 = _RAND_1078[7:0];
  _RAND_1079 = {1{`RANDOM}};
  lineBuffer_1072 = _RAND_1079[7:0];
  _RAND_1080 = {1{`RANDOM}};
  lineBuffer_1073 = _RAND_1080[7:0];
  _RAND_1081 = {1{`RANDOM}};
  lineBuffer_1074 = _RAND_1081[7:0];
  _RAND_1082 = {1{`RANDOM}};
  lineBuffer_1075 = _RAND_1082[7:0];
  _RAND_1083 = {1{`RANDOM}};
  lineBuffer_1076 = _RAND_1083[7:0];
  _RAND_1084 = {1{`RANDOM}};
  lineBuffer_1077 = _RAND_1084[7:0];
  _RAND_1085 = {1{`RANDOM}};
  lineBuffer_1078 = _RAND_1085[7:0];
  _RAND_1086 = {1{`RANDOM}};
  lineBuffer_1079 = _RAND_1086[7:0];
  _RAND_1087 = {1{`RANDOM}};
  lineBuffer_1080 = _RAND_1087[7:0];
  _RAND_1088 = {1{`RANDOM}};
  lineBuffer_1081 = _RAND_1088[7:0];
  _RAND_1089 = {1{`RANDOM}};
  lineBuffer_1082 = _RAND_1089[7:0];
  _RAND_1090 = {1{`RANDOM}};
  lineBuffer_1083 = _RAND_1090[7:0];
  _RAND_1091 = {1{`RANDOM}};
  lineBuffer_1084 = _RAND_1091[7:0];
  _RAND_1092 = {1{`RANDOM}};
  lineBuffer_1085 = _RAND_1092[7:0];
  _RAND_1093 = {1{`RANDOM}};
  lineBuffer_1086 = _RAND_1093[7:0];
  _RAND_1094 = {1{`RANDOM}};
  lineBuffer_1087 = _RAND_1094[7:0];
  _RAND_1095 = {1{`RANDOM}};
  lineBuffer_1088 = _RAND_1095[7:0];
  _RAND_1096 = {1{`RANDOM}};
  lineBuffer_1089 = _RAND_1096[7:0];
  _RAND_1097 = {1{`RANDOM}};
  lineBuffer_1090 = _RAND_1097[7:0];
  _RAND_1098 = {1{`RANDOM}};
  lineBuffer_1091 = _RAND_1098[7:0];
  _RAND_1099 = {1{`RANDOM}};
  lineBuffer_1092 = _RAND_1099[7:0];
  _RAND_1100 = {1{`RANDOM}};
  lineBuffer_1093 = _RAND_1100[7:0];
  _RAND_1101 = {1{`RANDOM}};
  lineBuffer_1094 = _RAND_1101[7:0];
  _RAND_1102 = {1{`RANDOM}};
  lineBuffer_1095 = _RAND_1102[7:0];
  _RAND_1103 = {1{`RANDOM}};
  lineBuffer_1096 = _RAND_1103[7:0];
  _RAND_1104 = {1{`RANDOM}};
  lineBuffer_1097 = _RAND_1104[7:0];
  _RAND_1105 = {1{`RANDOM}};
  lineBuffer_1098 = _RAND_1105[7:0];
  _RAND_1106 = {1{`RANDOM}};
  lineBuffer_1099 = _RAND_1106[7:0];
  _RAND_1107 = {1{`RANDOM}};
  lineBuffer_1100 = _RAND_1107[7:0];
  _RAND_1108 = {1{`RANDOM}};
  lineBuffer_1101 = _RAND_1108[7:0];
  _RAND_1109 = {1{`RANDOM}};
  lineBuffer_1102 = _RAND_1109[7:0];
  _RAND_1110 = {1{`RANDOM}};
  lineBuffer_1103 = _RAND_1110[7:0];
  _RAND_1111 = {1{`RANDOM}};
  lineBuffer_1104 = _RAND_1111[7:0];
  _RAND_1112 = {1{`RANDOM}};
  lineBuffer_1105 = _RAND_1112[7:0];
  _RAND_1113 = {1{`RANDOM}};
  lineBuffer_1106 = _RAND_1113[7:0];
  _RAND_1114 = {1{`RANDOM}};
  lineBuffer_1107 = _RAND_1114[7:0];
  _RAND_1115 = {1{`RANDOM}};
  lineBuffer_1108 = _RAND_1115[7:0];
  _RAND_1116 = {1{`RANDOM}};
  lineBuffer_1109 = _RAND_1116[7:0];
  _RAND_1117 = {1{`RANDOM}};
  lineBuffer_1110 = _RAND_1117[7:0];
  _RAND_1118 = {1{`RANDOM}};
  lineBuffer_1111 = _RAND_1118[7:0];
  _RAND_1119 = {1{`RANDOM}};
  lineBuffer_1112 = _RAND_1119[7:0];
  _RAND_1120 = {1{`RANDOM}};
  lineBuffer_1113 = _RAND_1120[7:0];
  _RAND_1121 = {1{`RANDOM}};
  lineBuffer_1114 = _RAND_1121[7:0];
  _RAND_1122 = {1{`RANDOM}};
  lineBuffer_1115 = _RAND_1122[7:0];
  _RAND_1123 = {1{`RANDOM}};
  lineBuffer_1116 = _RAND_1123[7:0];
  _RAND_1124 = {1{`RANDOM}};
  lineBuffer_1117 = _RAND_1124[7:0];
  _RAND_1125 = {1{`RANDOM}};
  lineBuffer_1118 = _RAND_1125[7:0];
  _RAND_1126 = {1{`RANDOM}};
  lineBuffer_1119 = _RAND_1126[7:0];
  _RAND_1127 = {1{`RANDOM}};
  lineBuffer_1120 = _RAND_1127[7:0];
  _RAND_1128 = {1{`RANDOM}};
  lineBuffer_1121 = _RAND_1128[7:0];
  _RAND_1129 = {1{`RANDOM}};
  lineBuffer_1122 = _RAND_1129[7:0];
  _RAND_1130 = {1{`RANDOM}};
  lineBuffer_1123 = _RAND_1130[7:0];
  _RAND_1131 = {1{`RANDOM}};
  lineBuffer_1124 = _RAND_1131[7:0];
  _RAND_1132 = {1{`RANDOM}};
  lineBuffer_1125 = _RAND_1132[7:0];
  _RAND_1133 = {1{`RANDOM}};
  lineBuffer_1126 = _RAND_1133[7:0];
  _RAND_1134 = {1{`RANDOM}};
  lineBuffer_1127 = _RAND_1134[7:0];
  _RAND_1135 = {1{`RANDOM}};
  lineBuffer_1128 = _RAND_1135[7:0];
  _RAND_1136 = {1{`RANDOM}};
  lineBuffer_1129 = _RAND_1136[7:0];
  _RAND_1137 = {1{`RANDOM}};
  lineBuffer_1130 = _RAND_1137[7:0];
  _RAND_1138 = {1{`RANDOM}};
  lineBuffer_1131 = _RAND_1138[7:0];
  _RAND_1139 = {1{`RANDOM}};
  lineBuffer_1132 = _RAND_1139[7:0];
  _RAND_1140 = {1{`RANDOM}};
  lineBuffer_1133 = _RAND_1140[7:0];
  _RAND_1141 = {1{`RANDOM}};
  lineBuffer_1134 = _RAND_1141[7:0];
  _RAND_1142 = {1{`RANDOM}};
  lineBuffer_1135 = _RAND_1142[7:0];
  _RAND_1143 = {1{`RANDOM}};
  lineBuffer_1136 = _RAND_1143[7:0];
  _RAND_1144 = {1{`RANDOM}};
  lineBuffer_1137 = _RAND_1144[7:0];
  _RAND_1145 = {1{`RANDOM}};
  lineBuffer_1138 = _RAND_1145[7:0];
  _RAND_1146 = {1{`RANDOM}};
  lineBuffer_1139 = _RAND_1146[7:0];
  _RAND_1147 = {1{`RANDOM}};
  lineBuffer_1140 = _RAND_1147[7:0];
  _RAND_1148 = {1{`RANDOM}};
  lineBuffer_1141 = _RAND_1148[7:0];
  _RAND_1149 = {1{`RANDOM}};
  lineBuffer_1142 = _RAND_1149[7:0];
  _RAND_1150 = {1{`RANDOM}};
  lineBuffer_1143 = _RAND_1150[7:0];
  _RAND_1151 = {1{`RANDOM}};
  lineBuffer_1144 = _RAND_1151[7:0];
  _RAND_1152 = {1{`RANDOM}};
  lineBuffer_1145 = _RAND_1152[7:0];
  _RAND_1153 = {1{`RANDOM}};
  lineBuffer_1146 = _RAND_1153[7:0];
  _RAND_1154 = {1{`RANDOM}};
  lineBuffer_1147 = _RAND_1154[7:0];
  _RAND_1155 = {1{`RANDOM}};
  lineBuffer_1148 = _RAND_1155[7:0];
  _RAND_1156 = {1{`RANDOM}};
  lineBuffer_1149 = _RAND_1156[7:0];
  _RAND_1157 = {1{`RANDOM}};
  lineBuffer_1150 = _RAND_1157[7:0];
  _RAND_1158 = {1{`RANDOM}};
  lineBuffer_1151 = _RAND_1158[7:0];
  _RAND_1159 = {1{`RANDOM}};
  lineBuffer_1152 = _RAND_1159[7:0];
  _RAND_1160 = {1{`RANDOM}};
  lineBuffer_1153 = _RAND_1160[7:0];
  _RAND_1161 = {1{`RANDOM}};
  lineBuffer_1154 = _RAND_1161[7:0];
  _RAND_1162 = {1{`RANDOM}};
  lineBuffer_1155 = _RAND_1162[7:0];
  _RAND_1163 = {1{`RANDOM}};
  lineBuffer_1156 = _RAND_1163[7:0];
  _RAND_1164 = {1{`RANDOM}};
  lineBuffer_1157 = _RAND_1164[7:0];
  _RAND_1165 = {1{`RANDOM}};
  lineBuffer_1158 = _RAND_1165[7:0];
  _RAND_1166 = {1{`RANDOM}};
  lineBuffer_1159 = _RAND_1166[7:0];
  _RAND_1167 = {1{`RANDOM}};
  lineBuffer_1160 = _RAND_1167[7:0];
  _RAND_1168 = {1{`RANDOM}};
  lineBuffer_1161 = _RAND_1168[7:0];
  _RAND_1169 = {1{`RANDOM}};
  lineBuffer_1162 = _RAND_1169[7:0];
  _RAND_1170 = {1{`RANDOM}};
  lineBuffer_1163 = _RAND_1170[7:0];
  _RAND_1171 = {1{`RANDOM}};
  lineBuffer_1164 = _RAND_1171[7:0];
  _RAND_1172 = {1{`RANDOM}};
  lineBuffer_1165 = _RAND_1172[7:0];
  _RAND_1173 = {1{`RANDOM}};
  lineBuffer_1166 = _RAND_1173[7:0];
  _RAND_1174 = {1{`RANDOM}};
  lineBuffer_1167 = _RAND_1174[7:0];
  _RAND_1175 = {1{`RANDOM}};
  lineBuffer_1168 = _RAND_1175[7:0];
  _RAND_1176 = {1{`RANDOM}};
  lineBuffer_1169 = _RAND_1176[7:0];
  _RAND_1177 = {1{`RANDOM}};
  lineBuffer_1170 = _RAND_1177[7:0];
  _RAND_1178 = {1{`RANDOM}};
  lineBuffer_1171 = _RAND_1178[7:0];
  _RAND_1179 = {1{`RANDOM}};
  lineBuffer_1172 = _RAND_1179[7:0];
  _RAND_1180 = {1{`RANDOM}};
  lineBuffer_1173 = _RAND_1180[7:0];
  _RAND_1181 = {1{`RANDOM}};
  lineBuffer_1174 = _RAND_1181[7:0];
  _RAND_1182 = {1{`RANDOM}};
  lineBuffer_1175 = _RAND_1182[7:0];
  _RAND_1183 = {1{`RANDOM}};
  lineBuffer_1176 = _RAND_1183[7:0];
  _RAND_1184 = {1{`RANDOM}};
  lineBuffer_1177 = _RAND_1184[7:0];
  _RAND_1185 = {1{`RANDOM}};
  lineBuffer_1178 = _RAND_1185[7:0];
  _RAND_1186 = {1{`RANDOM}};
  lineBuffer_1179 = _RAND_1186[7:0];
  _RAND_1187 = {1{`RANDOM}};
  lineBuffer_1180 = _RAND_1187[7:0];
  _RAND_1188 = {1{`RANDOM}};
  lineBuffer_1181 = _RAND_1188[7:0];
  _RAND_1189 = {1{`RANDOM}};
  lineBuffer_1182 = _RAND_1189[7:0];
  _RAND_1190 = {1{`RANDOM}};
  lineBuffer_1183 = _RAND_1190[7:0];
  _RAND_1191 = {1{`RANDOM}};
  lineBuffer_1184 = _RAND_1191[7:0];
  _RAND_1192 = {1{`RANDOM}};
  lineBuffer_1185 = _RAND_1192[7:0];
  _RAND_1193 = {1{`RANDOM}};
  lineBuffer_1186 = _RAND_1193[7:0];
  _RAND_1194 = {1{`RANDOM}};
  lineBuffer_1187 = _RAND_1194[7:0];
  _RAND_1195 = {1{`RANDOM}};
  lineBuffer_1188 = _RAND_1195[7:0];
  _RAND_1196 = {1{`RANDOM}};
  lineBuffer_1189 = _RAND_1196[7:0];
  _RAND_1197 = {1{`RANDOM}};
  lineBuffer_1190 = _RAND_1197[7:0];
  _RAND_1198 = {1{`RANDOM}};
  lineBuffer_1191 = _RAND_1198[7:0];
  _RAND_1199 = {1{`RANDOM}};
  lineBuffer_1192 = _RAND_1199[7:0];
  _RAND_1200 = {1{`RANDOM}};
  lineBuffer_1193 = _RAND_1200[7:0];
  _RAND_1201 = {1{`RANDOM}};
  lineBuffer_1194 = _RAND_1201[7:0];
  _RAND_1202 = {1{`RANDOM}};
  lineBuffer_1195 = _RAND_1202[7:0];
  _RAND_1203 = {1{`RANDOM}};
  lineBuffer_1196 = _RAND_1203[7:0];
  _RAND_1204 = {1{`RANDOM}};
  lineBuffer_1197 = _RAND_1204[7:0];
  _RAND_1205 = {1{`RANDOM}};
  lineBuffer_1198 = _RAND_1205[7:0];
  _RAND_1206 = {1{`RANDOM}};
  lineBuffer_1199 = _RAND_1206[7:0];
  _RAND_1207 = {1{`RANDOM}};
  lineBuffer_1200 = _RAND_1207[7:0];
  _RAND_1208 = {1{`RANDOM}};
  lineBuffer_1201 = _RAND_1208[7:0];
  _RAND_1209 = {1{`RANDOM}};
  lineBuffer_1202 = _RAND_1209[7:0];
  _RAND_1210 = {1{`RANDOM}};
  lineBuffer_1203 = _RAND_1210[7:0];
  _RAND_1211 = {1{`RANDOM}};
  lineBuffer_1204 = _RAND_1211[7:0];
  _RAND_1212 = {1{`RANDOM}};
  lineBuffer_1205 = _RAND_1212[7:0];
  _RAND_1213 = {1{`RANDOM}};
  lineBuffer_1206 = _RAND_1213[7:0];
  _RAND_1214 = {1{`RANDOM}};
  lineBuffer_1207 = _RAND_1214[7:0];
  _RAND_1215 = {1{`RANDOM}};
  lineBuffer_1208 = _RAND_1215[7:0];
  _RAND_1216 = {1{`RANDOM}};
  lineBuffer_1209 = _RAND_1216[7:0];
  _RAND_1217 = {1{`RANDOM}};
  lineBuffer_1210 = _RAND_1217[7:0];
  _RAND_1218 = {1{`RANDOM}};
  lineBuffer_1211 = _RAND_1218[7:0];
  _RAND_1219 = {1{`RANDOM}};
  lineBuffer_1212 = _RAND_1219[7:0];
  _RAND_1220 = {1{`RANDOM}};
  lineBuffer_1213 = _RAND_1220[7:0];
  _RAND_1221 = {1{`RANDOM}};
  lineBuffer_1214 = _RAND_1221[7:0];
  _RAND_1222 = {1{`RANDOM}};
  lineBuffer_1215 = _RAND_1222[7:0];
  _RAND_1223 = {1{`RANDOM}};
  lineBuffer_1216 = _RAND_1223[7:0];
  _RAND_1224 = {1{`RANDOM}};
  lineBuffer_1217 = _RAND_1224[7:0];
  _RAND_1225 = {1{`RANDOM}};
  lineBuffer_1218 = _RAND_1225[7:0];
  _RAND_1226 = {1{`RANDOM}};
  lineBuffer_1219 = _RAND_1226[7:0];
  _RAND_1227 = {1{`RANDOM}};
  lineBuffer_1220 = _RAND_1227[7:0];
  _RAND_1228 = {1{`RANDOM}};
  lineBuffer_1221 = _RAND_1228[7:0];
  _RAND_1229 = {1{`RANDOM}};
  lineBuffer_1222 = _RAND_1229[7:0];
  _RAND_1230 = {1{`RANDOM}};
  lineBuffer_1223 = _RAND_1230[7:0];
  _RAND_1231 = {1{`RANDOM}};
  lineBuffer_1224 = _RAND_1231[7:0];
  _RAND_1232 = {1{`RANDOM}};
  lineBuffer_1225 = _RAND_1232[7:0];
  _RAND_1233 = {1{`RANDOM}};
  lineBuffer_1226 = _RAND_1233[7:0];
  _RAND_1234 = {1{`RANDOM}};
  lineBuffer_1227 = _RAND_1234[7:0];
  _RAND_1235 = {1{`RANDOM}};
  lineBuffer_1228 = _RAND_1235[7:0];
  _RAND_1236 = {1{`RANDOM}};
  lineBuffer_1229 = _RAND_1236[7:0];
  _RAND_1237 = {1{`RANDOM}};
  lineBuffer_1230 = _RAND_1237[7:0];
  _RAND_1238 = {1{`RANDOM}};
  lineBuffer_1231 = _RAND_1238[7:0];
  _RAND_1239 = {1{`RANDOM}};
  lineBuffer_1232 = _RAND_1239[7:0];
  _RAND_1240 = {1{`RANDOM}};
  lineBuffer_1233 = _RAND_1240[7:0];
  _RAND_1241 = {1{`RANDOM}};
  lineBuffer_1234 = _RAND_1241[7:0];
  _RAND_1242 = {1{`RANDOM}};
  lineBuffer_1235 = _RAND_1242[7:0];
  _RAND_1243 = {1{`RANDOM}};
  lineBuffer_1236 = _RAND_1243[7:0];
  _RAND_1244 = {1{`RANDOM}};
  lineBuffer_1237 = _RAND_1244[7:0];
  _RAND_1245 = {1{`RANDOM}};
  lineBuffer_1238 = _RAND_1245[7:0];
  _RAND_1246 = {1{`RANDOM}};
  lineBuffer_1239 = _RAND_1246[7:0];
  _RAND_1247 = {1{`RANDOM}};
  lineBuffer_1240 = _RAND_1247[7:0];
  _RAND_1248 = {1{`RANDOM}};
  lineBuffer_1241 = _RAND_1248[7:0];
  _RAND_1249 = {1{`RANDOM}};
  lineBuffer_1242 = _RAND_1249[7:0];
  _RAND_1250 = {1{`RANDOM}};
  lineBuffer_1243 = _RAND_1250[7:0];
  _RAND_1251 = {1{`RANDOM}};
  lineBuffer_1244 = _RAND_1251[7:0];
  _RAND_1252 = {1{`RANDOM}};
  lineBuffer_1245 = _RAND_1252[7:0];
  _RAND_1253 = {1{`RANDOM}};
  lineBuffer_1246 = _RAND_1253[7:0];
  _RAND_1254 = {1{`RANDOM}};
  lineBuffer_1247 = _RAND_1254[7:0];
  _RAND_1255 = {1{`RANDOM}};
  lineBuffer_1248 = _RAND_1255[7:0];
  _RAND_1256 = {1{`RANDOM}};
  lineBuffer_1249 = _RAND_1256[7:0];
  _RAND_1257 = {1{`RANDOM}};
  lineBuffer_1250 = _RAND_1257[7:0];
  _RAND_1258 = {1{`RANDOM}};
  lineBuffer_1251 = _RAND_1258[7:0];
  _RAND_1259 = {1{`RANDOM}};
  lineBuffer_1252 = _RAND_1259[7:0];
  _RAND_1260 = {1{`RANDOM}};
  lineBuffer_1253 = _RAND_1260[7:0];
  _RAND_1261 = {1{`RANDOM}};
  lineBuffer_1254 = _RAND_1261[7:0];
  _RAND_1262 = {1{`RANDOM}};
  lineBuffer_1255 = _RAND_1262[7:0];
  _RAND_1263 = {1{`RANDOM}};
  lineBuffer_1256 = _RAND_1263[7:0];
  _RAND_1264 = {1{`RANDOM}};
  lineBuffer_1257 = _RAND_1264[7:0];
  _RAND_1265 = {1{`RANDOM}};
  lineBuffer_1258 = _RAND_1265[7:0];
  _RAND_1266 = {1{`RANDOM}};
  lineBuffer_1259 = _RAND_1266[7:0];
  _RAND_1267 = {1{`RANDOM}};
  lineBuffer_1260 = _RAND_1267[7:0];
  _RAND_1268 = {1{`RANDOM}};
  lineBuffer_1261 = _RAND_1268[7:0];
  _RAND_1269 = {1{`RANDOM}};
  lineBuffer_1262 = _RAND_1269[7:0];
  _RAND_1270 = {1{`RANDOM}};
  lineBuffer_1263 = _RAND_1270[7:0];
  _RAND_1271 = {1{`RANDOM}};
  lineBuffer_1264 = _RAND_1271[7:0];
  _RAND_1272 = {1{`RANDOM}};
  lineBuffer_1265 = _RAND_1272[7:0];
  _RAND_1273 = {1{`RANDOM}};
  lineBuffer_1266 = _RAND_1273[7:0];
  _RAND_1274 = {1{`RANDOM}};
  lineBuffer_1267 = _RAND_1274[7:0];
  _RAND_1275 = {1{`RANDOM}};
  lineBuffer_1268 = _RAND_1275[7:0];
  _RAND_1276 = {1{`RANDOM}};
  lineBuffer_1269 = _RAND_1276[7:0];
  _RAND_1277 = {1{`RANDOM}};
  lineBuffer_1270 = _RAND_1277[7:0];
  _RAND_1278 = {1{`RANDOM}};
  lineBuffer_1271 = _RAND_1278[7:0];
  _RAND_1279 = {1{`RANDOM}};
  lineBuffer_1272 = _RAND_1279[7:0];
  _RAND_1280 = {1{`RANDOM}};
  lineBuffer_1273 = _RAND_1280[7:0];
  _RAND_1281 = {1{`RANDOM}};
  lineBuffer_1274 = _RAND_1281[7:0];
  _RAND_1282 = {1{`RANDOM}};
  lineBuffer_1275 = _RAND_1282[7:0];
  _RAND_1283 = {1{`RANDOM}};
  lineBuffer_1276 = _RAND_1283[7:0];
  _RAND_1284 = {1{`RANDOM}};
  lineBuffer_1277 = _RAND_1284[7:0];
  _RAND_1285 = {1{`RANDOM}};
  lineBuffer_1278 = _RAND_1285[7:0];
  _RAND_1286 = {1{`RANDOM}};
  lineBuffer_1279 = _RAND_1286[7:0];
  _RAND_1287 = {1{`RANDOM}};
  lineBuffer_1280 = _RAND_1287[7:0];
  _RAND_1288 = {1{`RANDOM}};
  lineBuffer_1281 = _RAND_1288[7:0];
  _RAND_1289 = {1{`RANDOM}};
  lineBuffer_1282 = _RAND_1289[7:0];
  _RAND_1290 = {1{`RANDOM}};
  lineBuffer_1283 = _RAND_1290[7:0];
  _RAND_1291 = {1{`RANDOM}};
  lineBuffer_1284 = _RAND_1291[7:0];
  _RAND_1292 = {1{`RANDOM}};
  lineBuffer_1285 = _RAND_1292[7:0];
  _RAND_1293 = {1{`RANDOM}};
  lineBuffer_1286 = _RAND_1293[7:0];
  _RAND_1294 = {1{`RANDOM}};
  lineBuffer_1287 = _RAND_1294[7:0];
  _RAND_1295 = {1{`RANDOM}};
  lineBuffer_1288 = _RAND_1295[7:0];
  _RAND_1296 = {1{`RANDOM}};
  lineBuffer_1289 = _RAND_1296[7:0];
  _RAND_1297 = {1{`RANDOM}};
  lineBuffer_1290 = _RAND_1297[7:0];
  _RAND_1298 = {1{`RANDOM}};
  lineBuffer_1291 = _RAND_1298[7:0];
  _RAND_1299 = {1{`RANDOM}};
  lineBuffer_1292 = _RAND_1299[7:0];
  _RAND_1300 = {1{`RANDOM}};
  lineBuffer_1293 = _RAND_1300[7:0];
  _RAND_1301 = {1{`RANDOM}};
  lineBuffer_1294 = _RAND_1301[7:0];
  _RAND_1302 = {1{`RANDOM}};
  lineBuffer_1295 = _RAND_1302[7:0];
  _RAND_1303 = {1{`RANDOM}};
  lineBuffer_1296 = _RAND_1303[7:0];
  _RAND_1304 = {1{`RANDOM}};
  lineBuffer_1297 = _RAND_1304[7:0];
  _RAND_1305 = {1{`RANDOM}};
  lineBuffer_1298 = _RAND_1305[7:0];
  _RAND_1306 = {1{`RANDOM}};
  lineBuffer_1299 = _RAND_1306[7:0];
  _RAND_1307 = {1{`RANDOM}};
  lineBuffer_1300 = _RAND_1307[7:0];
  _RAND_1308 = {1{`RANDOM}};
  lineBuffer_1301 = _RAND_1308[7:0];
  _RAND_1309 = {1{`RANDOM}};
  lineBuffer_1302 = _RAND_1309[7:0];
  _RAND_1310 = {1{`RANDOM}};
  lineBuffer_1303 = _RAND_1310[7:0];
  _RAND_1311 = {1{`RANDOM}};
  lineBuffer_1304 = _RAND_1311[7:0];
  _RAND_1312 = {1{`RANDOM}};
  lineBuffer_1305 = _RAND_1312[7:0];
  _RAND_1313 = {1{`RANDOM}};
  lineBuffer_1306 = _RAND_1313[7:0];
  _RAND_1314 = {1{`RANDOM}};
  lineBuffer_1307 = _RAND_1314[7:0];
  _RAND_1315 = {1{`RANDOM}};
  lineBuffer_1308 = _RAND_1315[7:0];
  _RAND_1316 = {1{`RANDOM}};
  lineBuffer_1309 = _RAND_1316[7:0];
  _RAND_1317 = {1{`RANDOM}};
  lineBuffer_1310 = _RAND_1317[7:0];
  _RAND_1318 = {1{`RANDOM}};
  lineBuffer_1311 = _RAND_1318[7:0];
  _RAND_1319 = {1{`RANDOM}};
  lineBuffer_1312 = _RAND_1319[7:0];
  _RAND_1320 = {1{`RANDOM}};
  lineBuffer_1313 = _RAND_1320[7:0];
  _RAND_1321 = {1{`RANDOM}};
  lineBuffer_1314 = _RAND_1321[7:0];
  _RAND_1322 = {1{`RANDOM}};
  lineBuffer_1315 = _RAND_1322[7:0];
  _RAND_1323 = {1{`RANDOM}};
  lineBuffer_1316 = _RAND_1323[7:0];
  _RAND_1324 = {1{`RANDOM}};
  lineBuffer_1317 = _RAND_1324[7:0];
  _RAND_1325 = {1{`RANDOM}};
  lineBuffer_1318 = _RAND_1325[7:0];
  _RAND_1326 = {1{`RANDOM}};
  lineBuffer_1319 = _RAND_1326[7:0];
  _RAND_1327 = {1{`RANDOM}};
  lineBuffer_1320 = _RAND_1327[7:0];
  _RAND_1328 = {1{`RANDOM}};
  lineBuffer_1321 = _RAND_1328[7:0];
  _RAND_1329 = {1{`RANDOM}};
  lineBuffer_1322 = _RAND_1329[7:0];
  _RAND_1330 = {1{`RANDOM}};
  lineBuffer_1323 = _RAND_1330[7:0];
  _RAND_1331 = {1{`RANDOM}};
  lineBuffer_1324 = _RAND_1331[7:0];
  _RAND_1332 = {1{`RANDOM}};
  lineBuffer_1325 = _RAND_1332[7:0];
  _RAND_1333 = {1{`RANDOM}};
  lineBuffer_1326 = _RAND_1333[7:0];
  _RAND_1334 = {1{`RANDOM}};
  lineBuffer_1327 = _RAND_1334[7:0];
  _RAND_1335 = {1{`RANDOM}};
  lineBuffer_1328 = _RAND_1335[7:0];
  _RAND_1336 = {1{`RANDOM}};
  lineBuffer_1329 = _RAND_1336[7:0];
  _RAND_1337 = {1{`RANDOM}};
  lineBuffer_1330 = _RAND_1337[7:0];
  _RAND_1338 = {1{`RANDOM}};
  lineBuffer_1331 = _RAND_1338[7:0];
  _RAND_1339 = {1{`RANDOM}};
  lineBuffer_1332 = _RAND_1339[7:0];
  _RAND_1340 = {1{`RANDOM}};
  lineBuffer_1333 = _RAND_1340[7:0];
  _RAND_1341 = {1{`RANDOM}};
  lineBuffer_1334 = _RAND_1341[7:0];
  _RAND_1342 = {1{`RANDOM}};
  lineBuffer_1335 = _RAND_1342[7:0];
  _RAND_1343 = {1{`RANDOM}};
  lineBuffer_1336 = _RAND_1343[7:0];
  _RAND_1344 = {1{`RANDOM}};
  lineBuffer_1337 = _RAND_1344[7:0];
  _RAND_1345 = {1{`RANDOM}};
  lineBuffer_1338 = _RAND_1345[7:0];
  _RAND_1346 = {1{`RANDOM}};
  lineBuffer_1339 = _RAND_1346[7:0];
  _RAND_1347 = {1{`RANDOM}};
  lineBuffer_1340 = _RAND_1347[7:0];
  _RAND_1348 = {1{`RANDOM}};
  lineBuffer_1341 = _RAND_1348[7:0];
  _RAND_1349 = {1{`RANDOM}};
  lineBuffer_1342 = _RAND_1349[7:0];
  _RAND_1350 = {1{`RANDOM}};
  lineBuffer_1343 = _RAND_1350[7:0];
  _RAND_1351 = {1{`RANDOM}};
  lineBuffer_1344 = _RAND_1351[7:0];
  _RAND_1352 = {1{`RANDOM}};
  lineBuffer_1345 = _RAND_1352[7:0];
  _RAND_1353 = {1{`RANDOM}};
  lineBuffer_1346 = _RAND_1353[7:0];
  _RAND_1354 = {1{`RANDOM}};
  lineBuffer_1347 = _RAND_1354[7:0];
  _RAND_1355 = {1{`RANDOM}};
  lineBuffer_1348 = _RAND_1355[7:0];
  _RAND_1356 = {1{`RANDOM}};
  lineBuffer_1349 = _RAND_1356[7:0];
  _RAND_1357 = {1{`RANDOM}};
  lineBuffer_1350 = _RAND_1357[7:0];
  _RAND_1358 = {1{`RANDOM}};
  lineBuffer_1351 = _RAND_1358[7:0];
  _RAND_1359 = {1{`RANDOM}};
  lineBuffer_1352 = _RAND_1359[7:0];
  _RAND_1360 = {1{`RANDOM}};
  lineBuffer_1353 = _RAND_1360[7:0];
  _RAND_1361 = {1{`RANDOM}};
  lineBuffer_1354 = _RAND_1361[7:0];
  _RAND_1362 = {1{`RANDOM}};
  lineBuffer_1355 = _RAND_1362[7:0];
  _RAND_1363 = {1{`RANDOM}};
  lineBuffer_1356 = _RAND_1363[7:0];
  _RAND_1364 = {1{`RANDOM}};
  lineBuffer_1357 = _RAND_1364[7:0];
  _RAND_1365 = {1{`RANDOM}};
  lineBuffer_1358 = _RAND_1365[7:0];
  _RAND_1366 = {1{`RANDOM}};
  lineBuffer_1359 = _RAND_1366[7:0];
  _RAND_1367 = {1{`RANDOM}};
  lineBuffer_1360 = _RAND_1367[7:0];
  _RAND_1368 = {1{`RANDOM}};
  lineBuffer_1361 = _RAND_1368[7:0];
  _RAND_1369 = {1{`RANDOM}};
  lineBuffer_1362 = _RAND_1369[7:0];
  _RAND_1370 = {1{`RANDOM}};
  lineBuffer_1363 = _RAND_1370[7:0];
  _RAND_1371 = {1{`RANDOM}};
  lineBuffer_1364 = _RAND_1371[7:0];
  _RAND_1372 = {1{`RANDOM}};
  lineBuffer_1365 = _RAND_1372[7:0];
  _RAND_1373 = {1{`RANDOM}};
  lineBuffer_1366 = _RAND_1373[7:0];
  _RAND_1374 = {1{`RANDOM}};
  lineBuffer_1367 = _RAND_1374[7:0];
  _RAND_1375 = {1{`RANDOM}};
  lineBuffer_1368 = _RAND_1375[7:0];
  _RAND_1376 = {1{`RANDOM}};
  lineBuffer_1369 = _RAND_1376[7:0];
  _RAND_1377 = {1{`RANDOM}};
  lineBuffer_1370 = _RAND_1377[7:0];
  _RAND_1378 = {1{`RANDOM}};
  lineBuffer_1371 = _RAND_1378[7:0];
  _RAND_1379 = {1{`RANDOM}};
  lineBuffer_1372 = _RAND_1379[7:0];
  _RAND_1380 = {1{`RANDOM}};
  lineBuffer_1373 = _RAND_1380[7:0];
  _RAND_1381 = {1{`RANDOM}};
  lineBuffer_1374 = _RAND_1381[7:0];
  _RAND_1382 = {1{`RANDOM}};
  lineBuffer_1375 = _RAND_1382[7:0];
  _RAND_1383 = {1{`RANDOM}};
  lineBuffer_1376 = _RAND_1383[7:0];
  _RAND_1384 = {1{`RANDOM}};
  lineBuffer_1377 = _RAND_1384[7:0];
  _RAND_1385 = {1{`RANDOM}};
  lineBuffer_1378 = _RAND_1385[7:0];
  _RAND_1386 = {1{`RANDOM}};
  lineBuffer_1379 = _RAND_1386[7:0];
  _RAND_1387 = {1{`RANDOM}};
  lineBuffer_1380 = _RAND_1387[7:0];
  _RAND_1388 = {1{`RANDOM}};
  lineBuffer_1381 = _RAND_1388[7:0];
  _RAND_1389 = {1{`RANDOM}};
  lineBuffer_1382 = _RAND_1389[7:0];
  _RAND_1390 = {1{`RANDOM}};
  lineBuffer_1383 = _RAND_1390[7:0];
  _RAND_1391 = {1{`RANDOM}};
  lineBuffer_1384 = _RAND_1391[7:0];
  _RAND_1392 = {1{`RANDOM}};
  lineBuffer_1385 = _RAND_1392[7:0];
  _RAND_1393 = {1{`RANDOM}};
  lineBuffer_1386 = _RAND_1393[7:0];
  _RAND_1394 = {1{`RANDOM}};
  lineBuffer_1387 = _RAND_1394[7:0];
  _RAND_1395 = {1{`RANDOM}};
  lineBuffer_1388 = _RAND_1395[7:0];
  _RAND_1396 = {1{`RANDOM}};
  lineBuffer_1389 = _RAND_1396[7:0];
  _RAND_1397 = {1{`RANDOM}};
  lineBuffer_1390 = _RAND_1397[7:0];
  _RAND_1398 = {1{`RANDOM}};
  lineBuffer_1391 = _RAND_1398[7:0];
  _RAND_1399 = {1{`RANDOM}};
  lineBuffer_1392 = _RAND_1399[7:0];
  _RAND_1400 = {1{`RANDOM}};
  lineBuffer_1393 = _RAND_1400[7:0];
  _RAND_1401 = {1{`RANDOM}};
  lineBuffer_1394 = _RAND_1401[7:0];
  _RAND_1402 = {1{`RANDOM}};
  lineBuffer_1395 = _RAND_1402[7:0];
  _RAND_1403 = {1{`RANDOM}};
  lineBuffer_1396 = _RAND_1403[7:0];
  _RAND_1404 = {1{`RANDOM}};
  lineBuffer_1397 = _RAND_1404[7:0];
  _RAND_1405 = {1{`RANDOM}};
  lineBuffer_1398 = _RAND_1405[7:0];
  _RAND_1406 = {1{`RANDOM}};
  lineBuffer_1399 = _RAND_1406[7:0];
  _RAND_1407 = {1{`RANDOM}};
  lineBuffer_1400 = _RAND_1407[7:0];
  _RAND_1408 = {1{`RANDOM}};
  lineBuffer_1401 = _RAND_1408[7:0];
  _RAND_1409 = {1{`RANDOM}};
  lineBuffer_1402 = _RAND_1409[7:0];
  _RAND_1410 = {1{`RANDOM}};
  lineBuffer_1403 = _RAND_1410[7:0];
  _RAND_1411 = {1{`RANDOM}};
  lineBuffer_1404 = _RAND_1411[7:0];
  _RAND_1412 = {1{`RANDOM}};
  lineBuffer_1405 = _RAND_1412[7:0];
  _RAND_1413 = {1{`RANDOM}};
  lineBuffer_1406 = _RAND_1413[7:0];
  _RAND_1414 = {1{`RANDOM}};
  lineBuffer_1407 = _RAND_1414[7:0];
  _RAND_1415 = {1{`RANDOM}};
  lineBuffer_1408 = _RAND_1415[7:0];
  _RAND_1416 = {1{`RANDOM}};
  lineBuffer_1409 = _RAND_1416[7:0];
  _RAND_1417 = {1{`RANDOM}};
  lineBuffer_1410 = _RAND_1417[7:0];
  _RAND_1418 = {1{`RANDOM}};
  lineBuffer_1411 = _RAND_1418[7:0];
  _RAND_1419 = {1{`RANDOM}};
  lineBuffer_1412 = _RAND_1419[7:0];
  _RAND_1420 = {1{`RANDOM}};
  lineBuffer_1413 = _RAND_1420[7:0];
  _RAND_1421 = {1{`RANDOM}};
  lineBuffer_1414 = _RAND_1421[7:0];
  _RAND_1422 = {1{`RANDOM}};
  lineBuffer_1415 = _RAND_1422[7:0];
  _RAND_1423 = {1{`RANDOM}};
  lineBuffer_1416 = _RAND_1423[7:0];
  _RAND_1424 = {1{`RANDOM}};
  lineBuffer_1417 = _RAND_1424[7:0];
  _RAND_1425 = {1{`RANDOM}};
  lineBuffer_1418 = _RAND_1425[7:0];
  _RAND_1426 = {1{`RANDOM}};
  lineBuffer_1419 = _RAND_1426[7:0];
  _RAND_1427 = {1{`RANDOM}};
  lineBuffer_1420 = _RAND_1427[7:0];
  _RAND_1428 = {1{`RANDOM}};
  lineBuffer_1421 = _RAND_1428[7:0];
  _RAND_1429 = {1{`RANDOM}};
  lineBuffer_1422 = _RAND_1429[7:0];
  _RAND_1430 = {1{`RANDOM}};
  lineBuffer_1423 = _RAND_1430[7:0];
  _RAND_1431 = {1{`RANDOM}};
  lineBuffer_1424 = _RAND_1431[7:0];
  _RAND_1432 = {1{`RANDOM}};
  lineBuffer_1425 = _RAND_1432[7:0];
  _RAND_1433 = {1{`RANDOM}};
  lineBuffer_1426 = _RAND_1433[7:0];
  _RAND_1434 = {1{`RANDOM}};
  lineBuffer_1427 = _RAND_1434[7:0];
  _RAND_1435 = {1{`RANDOM}};
  lineBuffer_1428 = _RAND_1435[7:0];
  _RAND_1436 = {1{`RANDOM}};
  lineBuffer_1429 = _RAND_1436[7:0];
  _RAND_1437 = {1{`RANDOM}};
  lineBuffer_1430 = _RAND_1437[7:0];
  _RAND_1438 = {1{`RANDOM}};
  lineBuffer_1431 = _RAND_1438[7:0];
  _RAND_1439 = {1{`RANDOM}};
  lineBuffer_1432 = _RAND_1439[7:0];
  _RAND_1440 = {1{`RANDOM}};
  lineBuffer_1433 = _RAND_1440[7:0];
  _RAND_1441 = {1{`RANDOM}};
  lineBuffer_1434 = _RAND_1441[7:0];
  _RAND_1442 = {1{`RANDOM}};
  lineBuffer_1435 = _RAND_1442[7:0];
  _RAND_1443 = {1{`RANDOM}};
  lineBuffer_1436 = _RAND_1443[7:0];
  _RAND_1444 = {1{`RANDOM}};
  lineBuffer_1437 = _RAND_1444[7:0];
  _RAND_1445 = {1{`RANDOM}};
  lineBuffer_1438 = _RAND_1445[7:0];
  _RAND_1446 = {1{`RANDOM}};
  lineBuffer_1439 = _RAND_1446[7:0];
  _RAND_1447 = {1{`RANDOM}};
  lineBuffer_1440 = _RAND_1447[7:0];
  _RAND_1448 = {1{`RANDOM}};
  lineBuffer_1441 = _RAND_1448[7:0];
  _RAND_1449 = {1{`RANDOM}};
  lineBuffer_1442 = _RAND_1449[7:0];
  _RAND_1450 = {1{`RANDOM}};
  lineBuffer_1443 = _RAND_1450[7:0];
  _RAND_1451 = {1{`RANDOM}};
  lineBuffer_1444 = _RAND_1451[7:0];
  _RAND_1452 = {1{`RANDOM}};
  lineBuffer_1445 = _RAND_1452[7:0];
  _RAND_1453 = {1{`RANDOM}};
  lineBuffer_1446 = _RAND_1453[7:0];
  _RAND_1454 = {1{`RANDOM}};
  lineBuffer_1447 = _RAND_1454[7:0];
  _RAND_1455 = {1{`RANDOM}};
  lineBuffer_1448 = _RAND_1455[7:0];
  _RAND_1456 = {1{`RANDOM}};
  lineBuffer_1449 = _RAND_1456[7:0];
  _RAND_1457 = {1{`RANDOM}};
  lineBuffer_1450 = _RAND_1457[7:0];
  _RAND_1458 = {1{`RANDOM}};
  lineBuffer_1451 = _RAND_1458[7:0];
  _RAND_1459 = {1{`RANDOM}};
  lineBuffer_1452 = _RAND_1459[7:0];
  _RAND_1460 = {1{`RANDOM}};
  lineBuffer_1453 = _RAND_1460[7:0];
  _RAND_1461 = {1{`RANDOM}};
  lineBuffer_1454 = _RAND_1461[7:0];
  _RAND_1462 = {1{`RANDOM}};
  lineBuffer_1455 = _RAND_1462[7:0];
  _RAND_1463 = {1{`RANDOM}};
  lineBuffer_1456 = _RAND_1463[7:0];
  _RAND_1464 = {1{`RANDOM}};
  lineBuffer_1457 = _RAND_1464[7:0];
  _RAND_1465 = {1{`RANDOM}};
  lineBuffer_1458 = _RAND_1465[7:0];
  _RAND_1466 = {1{`RANDOM}};
  lineBuffer_1459 = _RAND_1466[7:0];
  _RAND_1467 = {1{`RANDOM}};
  lineBuffer_1460 = _RAND_1467[7:0];
  _RAND_1468 = {1{`RANDOM}};
  lineBuffer_1461 = _RAND_1468[7:0];
  _RAND_1469 = {1{`RANDOM}};
  lineBuffer_1462 = _RAND_1469[7:0];
  _RAND_1470 = {1{`RANDOM}};
  lineBuffer_1463 = _RAND_1470[7:0];
  _RAND_1471 = {1{`RANDOM}};
  lineBuffer_1464 = _RAND_1471[7:0];
  _RAND_1472 = {1{`RANDOM}};
  lineBuffer_1465 = _RAND_1472[7:0];
  _RAND_1473 = {1{`RANDOM}};
  lineBuffer_1466 = _RAND_1473[7:0];
  _RAND_1474 = {1{`RANDOM}};
  lineBuffer_1467 = _RAND_1474[7:0];
  _RAND_1475 = {1{`RANDOM}};
  lineBuffer_1468 = _RAND_1475[7:0];
  _RAND_1476 = {1{`RANDOM}};
  lineBuffer_1469 = _RAND_1476[7:0];
  _RAND_1477 = {1{`RANDOM}};
  lineBuffer_1470 = _RAND_1477[7:0];
  _RAND_1478 = {1{`RANDOM}};
  lineBuffer_1471 = _RAND_1478[7:0];
  _RAND_1479 = {1{`RANDOM}};
  lineBuffer_1472 = _RAND_1479[7:0];
  _RAND_1480 = {1{`RANDOM}};
  lineBuffer_1473 = _RAND_1480[7:0];
  _RAND_1481 = {1{`RANDOM}};
  lineBuffer_1474 = _RAND_1481[7:0];
  _RAND_1482 = {1{`RANDOM}};
  lineBuffer_1475 = _RAND_1482[7:0];
  _RAND_1483 = {1{`RANDOM}};
  lineBuffer_1476 = _RAND_1483[7:0];
  _RAND_1484 = {1{`RANDOM}};
  lineBuffer_1477 = _RAND_1484[7:0];
  _RAND_1485 = {1{`RANDOM}};
  lineBuffer_1478 = _RAND_1485[7:0];
  _RAND_1486 = {1{`RANDOM}};
  lineBuffer_1479 = _RAND_1486[7:0];
  _RAND_1487 = {1{`RANDOM}};
  lineBuffer_1480 = _RAND_1487[7:0];
  _RAND_1488 = {1{`RANDOM}};
  lineBuffer_1481 = _RAND_1488[7:0];
  _RAND_1489 = {1{`RANDOM}};
  lineBuffer_1482 = _RAND_1489[7:0];
  _RAND_1490 = {1{`RANDOM}};
  lineBuffer_1483 = _RAND_1490[7:0];
  _RAND_1491 = {1{`RANDOM}};
  lineBuffer_1484 = _RAND_1491[7:0];
  _RAND_1492 = {1{`RANDOM}};
  lineBuffer_1485 = _RAND_1492[7:0];
  _RAND_1493 = {1{`RANDOM}};
  lineBuffer_1486 = _RAND_1493[7:0];
  _RAND_1494 = {1{`RANDOM}};
  lineBuffer_1487 = _RAND_1494[7:0];
  _RAND_1495 = {1{`RANDOM}};
  lineBuffer_1488 = _RAND_1495[7:0];
  _RAND_1496 = {1{`RANDOM}};
  lineBuffer_1489 = _RAND_1496[7:0];
  _RAND_1497 = {1{`RANDOM}};
  lineBuffer_1490 = _RAND_1497[7:0];
  _RAND_1498 = {1{`RANDOM}};
  lineBuffer_1491 = _RAND_1498[7:0];
  _RAND_1499 = {1{`RANDOM}};
  lineBuffer_1492 = _RAND_1499[7:0];
  _RAND_1500 = {1{`RANDOM}};
  lineBuffer_1493 = _RAND_1500[7:0];
  _RAND_1501 = {1{`RANDOM}};
  lineBuffer_1494 = _RAND_1501[7:0];
  _RAND_1502 = {1{`RANDOM}};
  lineBuffer_1495 = _RAND_1502[7:0];
  _RAND_1503 = {1{`RANDOM}};
  lineBuffer_1496 = _RAND_1503[7:0];
  _RAND_1504 = {1{`RANDOM}};
  lineBuffer_1497 = _RAND_1504[7:0];
  _RAND_1505 = {1{`RANDOM}};
  lineBuffer_1498 = _RAND_1505[7:0];
  _RAND_1506 = {1{`RANDOM}};
  lineBuffer_1499 = _RAND_1506[7:0];
  _RAND_1507 = {1{`RANDOM}};
  lineBuffer_1500 = _RAND_1507[7:0];
  _RAND_1508 = {1{`RANDOM}};
  lineBuffer_1501 = _RAND_1508[7:0];
  _RAND_1509 = {1{`RANDOM}};
  lineBuffer_1502 = _RAND_1509[7:0];
  _RAND_1510 = {1{`RANDOM}};
  lineBuffer_1503 = _RAND_1510[7:0];
  _RAND_1511 = {1{`RANDOM}};
  lineBuffer_1504 = _RAND_1511[7:0];
  _RAND_1512 = {1{`RANDOM}};
  lineBuffer_1505 = _RAND_1512[7:0];
  _RAND_1513 = {1{`RANDOM}};
  lineBuffer_1506 = _RAND_1513[7:0];
  _RAND_1514 = {1{`RANDOM}};
  lineBuffer_1507 = _RAND_1514[7:0];
  _RAND_1515 = {1{`RANDOM}};
  lineBuffer_1508 = _RAND_1515[7:0];
  _RAND_1516 = {1{`RANDOM}};
  lineBuffer_1509 = _RAND_1516[7:0];
  _RAND_1517 = {1{`RANDOM}};
  lineBuffer_1510 = _RAND_1517[7:0];
  _RAND_1518 = {1{`RANDOM}};
  lineBuffer_1511 = _RAND_1518[7:0];
  _RAND_1519 = {1{`RANDOM}};
  lineBuffer_1512 = _RAND_1519[7:0];
  _RAND_1520 = {1{`RANDOM}};
  lineBuffer_1513 = _RAND_1520[7:0];
  _RAND_1521 = {1{`RANDOM}};
  lineBuffer_1514 = _RAND_1521[7:0];
  _RAND_1522 = {1{`RANDOM}};
  lineBuffer_1515 = _RAND_1522[7:0];
  _RAND_1523 = {1{`RANDOM}};
  lineBuffer_1516 = _RAND_1523[7:0];
  _RAND_1524 = {1{`RANDOM}};
  lineBuffer_1517 = _RAND_1524[7:0];
  _RAND_1525 = {1{`RANDOM}};
  lineBuffer_1518 = _RAND_1525[7:0];
  _RAND_1526 = {1{`RANDOM}};
  lineBuffer_1519 = _RAND_1526[7:0];
  _RAND_1527 = {1{`RANDOM}};
  lineBuffer_1520 = _RAND_1527[7:0];
  _RAND_1528 = {1{`RANDOM}};
  lineBuffer_1521 = _RAND_1528[7:0];
  _RAND_1529 = {1{`RANDOM}};
  lineBuffer_1522 = _RAND_1529[7:0];
  _RAND_1530 = {1{`RANDOM}};
  lineBuffer_1523 = _RAND_1530[7:0];
  _RAND_1531 = {1{`RANDOM}};
  lineBuffer_1524 = _RAND_1531[7:0];
  _RAND_1532 = {1{`RANDOM}};
  lineBuffer_1525 = _RAND_1532[7:0];
  _RAND_1533 = {1{`RANDOM}};
  lineBuffer_1526 = _RAND_1533[7:0];
  _RAND_1534 = {1{`RANDOM}};
  lineBuffer_1527 = _RAND_1534[7:0];
  _RAND_1535 = {1{`RANDOM}};
  lineBuffer_1528 = _RAND_1535[7:0];
  _RAND_1536 = {1{`RANDOM}};
  lineBuffer_1529 = _RAND_1536[7:0];
  _RAND_1537 = {1{`RANDOM}};
  lineBuffer_1530 = _RAND_1537[7:0];
  _RAND_1538 = {1{`RANDOM}};
  lineBuffer_1531 = _RAND_1538[7:0];
  _RAND_1539 = {1{`RANDOM}};
  lineBuffer_1532 = _RAND_1539[7:0];
  _RAND_1540 = {1{`RANDOM}};
  lineBuffer_1533 = _RAND_1540[7:0];
  _RAND_1541 = {1{`RANDOM}};
  lineBuffer_1534 = _RAND_1541[7:0];
  _RAND_1542 = {1{`RANDOM}};
  lineBuffer_1535 = _RAND_1542[7:0];
  _RAND_1543 = {1{`RANDOM}};
  lineBuffer_1536 = _RAND_1543[7:0];
  _RAND_1544 = {1{`RANDOM}};
  lineBuffer_1537 = _RAND_1544[7:0];
  _RAND_1545 = {1{`RANDOM}};
  lineBuffer_1538 = _RAND_1545[7:0];
  _RAND_1546 = {1{`RANDOM}};
  lineBuffer_1539 = _RAND_1546[7:0];
  _RAND_1547 = {1{`RANDOM}};
  lineBuffer_1540 = _RAND_1547[7:0];
  _RAND_1548 = {1{`RANDOM}};
  lineBuffer_1541 = _RAND_1548[7:0];
  _RAND_1549 = {1{`RANDOM}};
  lineBuffer_1542 = _RAND_1549[7:0];
  _RAND_1550 = {1{`RANDOM}};
  lineBuffer_1543 = _RAND_1550[7:0];
  _RAND_1551 = {1{`RANDOM}};
  lineBuffer_1544 = _RAND_1551[7:0];
  _RAND_1552 = {1{`RANDOM}};
  lineBuffer_1545 = _RAND_1552[7:0];
  _RAND_1553 = {1{`RANDOM}};
  lineBuffer_1546 = _RAND_1553[7:0];
  _RAND_1554 = {1{`RANDOM}};
  lineBuffer_1547 = _RAND_1554[7:0];
  _RAND_1555 = {1{`RANDOM}};
  lineBuffer_1548 = _RAND_1555[7:0];
  _RAND_1556 = {1{`RANDOM}};
  lineBuffer_1549 = _RAND_1556[7:0];
  _RAND_1557 = {1{`RANDOM}};
  lineBuffer_1550 = _RAND_1557[7:0];
  _RAND_1558 = {1{`RANDOM}};
  lineBuffer_1551 = _RAND_1558[7:0];
  _RAND_1559 = {1{`RANDOM}};
  lineBuffer_1552 = _RAND_1559[7:0];
  _RAND_1560 = {1{`RANDOM}};
  lineBuffer_1553 = _RAND_1560[7:0];
  _RAND_1561 = {1{`RANDOM}};
  lineBuffer_1554 = _RAND_1561[7:0];
  _RAND_1562 = {1{`RANDOM}};
  lineBuffer_1555 = _RAND_1562[7:0];
  _RAND_1563 = {1{`RANDOM}};
  lineBuffer_1556 = _RAND_1563[7:0];
  _RAND_1564 = {1{`RANDOM}};
  lineBuffer_1557 = _RAND_1564[7:0];
  _RAND_1565 = {1{`RANDOM}};
  lineBuffer_1558 = _RAND_1565[7:0];
  _RAND_1566 = {1{`RANDOM}};
  lineBuffer_1559 = _RAND_1566[7:0];
  _RAND_1567 = {1{`RANDOM}};
  lineBuffer_1560 = _RAND_1567[7:0];
  _RAND_1568 = {1{`RANDOM}};
  lineBuffer_1561 = _RAND_1568[7:0];
  _RAND_1569 = {1{`RANDOM}};
  lineBuffer_1562 = _RAND_1569[7:0];
  _RAND_1570 = {1{`RANDOM}};
  lineBuffer_1563 = _RAND_1570[7:0];
  _RAND_1571 = {1{`RANDOM}};
  lineBuffer_1564 = _RAND_1571[7:0];
  _RAND_1572 = {1{`RANDOM}};
  lineBuffer_1565 = _RAND_1572[7:0];
  _RAND_1573 = {1{`RANDOM}};
  lineBuffer_1566 = _RAND_1573[7:0];
  _RAND_1574 = {1{`RANDOM}};
  lineBuffer_1567 = _RAND_1574[7:0];
  _RAND_1575 = {1{`RANDOM}};
  lineBuffer_1568 = _RAND_1575[7:0];
  _RAND_1576 = {1{`RANDOM}};
  lineBuffer_1569 = _RAND_1576[7:0];
  _RAND_1577 = {1{`RANDOM}};
  lineBuffer_1570 = _RAND_1577[7:0];
  _RAND_1578 = {1{`RANDOM}};
  lineBuffer_1571 = _RAND_1578[7:0];
  _RAND_1579 = {1{`RANDOM}};
  lineBuffer_1572 = _RAND_1579[7:0];
  _RAND_1580 = {1{`RANDOM}};
  lineBuffer_1573 = _RAND_1580[7:0];
  _RAND_1581 = {1{`RANDOM}};
  lineBuffer_1574 = _RAND_1581[7:0];
  _RAND_1582 = {1{`RANDOM}};
  lineBuffer_1575 = _RAND_1582[7:0];
  _RAND_1583 = {1{`RANDOM}};
  lineBuffer_1576 = _RAND_1583[7:0];
  _RAND_1584 = {1{`RANDOM}};
  lineBuffer_1577 = _RAND_1584[7:0];
  _RAND_1585 = {1{`RANDOM}};
  lineBuffer_1578 = _RAND_1585[7:0];
  _RAND_1586 = {1{`RANDOM}};
  lineBuffer_1579 = _RAND_1586[7:0];
  _RAND_1587 = {1{`RANDOM}};
  lineBuffer_1580 = _RAND_1587[7:0];
  _RAND_1588 = {1{`RANDOM}};
  lineBuffer_1581 = _RAND_1588[7:0];
  _RAND_1589 = {1{`RANDOM}};
  lineBuffer_1582 = _RAND_1589[7:0];
  _RAND_1590 = {1{`RANDOM}};
  lineBuffer_1583 = _RAND_1590[7:0];
  _RAND_1591 = {1{`RANDOM}};
  lineBuffer_1584 = _RAND_1591[7:0];
  _RAND_1592 = {1{`RANDOM}};
  lineBuffer_1585 = _RAND_1592[7:0];
  _RAND_1593 = {1{`RANDOM}};
  lineBuffer_1586 = _RAND_1593[7:0];
  _RAND_1594 = {1{`RANDOM}};
  lineBuffer_1587 = _RAND_1594[7:0];
  _RAND_1595 = {1{`RANDOM}};
  lineBuffer_1588 = _RAND_1595[7:0];
  _RAND_1596 = {1{`RANDOM}};
  lineBuffer_1589 = _RAND_1596[7:0];
  _RAND_1597 = {1{`RANDOM}};
  lineBuffer_1590 = _RAND_1597[7:0];
  _RAND_1598 = {1{`RANDOM}};
  lineBuffer_1591 = _RAND_1598[7:0];
  _RAND_1599 = {1{`RANDOM}};
  lineBuffer_1592 = _RAND_1599[7:0];
  _RAND_1600 = {1{`RANDOM}};
  lineBuffer_1593 = _RAND_1600[7:0];
  _RAND_1601 = {1{`RANDOM}};
  lineBuffer_1594 = _RAND_1601[7:0];
  _RAND_1602 = {1{`RANDOM}};
  lineBuffer_1595 = _RAND_1602[7:0];
  _RAND_1603 = {1{`RANDOM}};
  lineBuffer_1596 = _RAND_1603[7:0];
  _RAND_1604 = {1{`RANDOM}};
  lineBuffer_1597 = _RAND_1604[7:0];
  _RAND_1605 = {1{`RANDOM}};
  lineBuffer_1598 = _RAND_1605[7:0];
  _RAND_1606 = {1{`RANDOM}};
  lineBuffer_1599 = _RAND_1606[7:0];
  _RAND_1607 = {1{`RANDOM}};
  lineBuffer_1600 = _RAND_1607[7:0];
  _RAND_1608 = {1{`RANDOM}};
  lineBuffer_1601 = _RAND_1608[7:0];
  _RAND_1609 = {1{`RANDOM}};
  lineBuffer_1602 = _RAND_1609[7:0];
  _RAND_1610 = {1{`RANDOM}};
  lineBuffer_1603 = _RAND_1610[7:0];
  _RAND_1611 = {1{`RANDOM}};
  lineBuffer_1604 = _RAND_1611[7:0];
  _RAND_1612 = {1{`RANDOM}};
  lineBuffer_1605 = _RAND_1612[7:0];
  _RAND_1613 = {1{`RANDOM}};
  lineBuffer_1606 = _RAND_1613[7:0];
  _RAND_1614 = {1{`RANDOM}};
  lineBuffer_1607 = _RAND_1614[7:0];
  _RAND_1615 = {1{`RANDOM}};
  lineBuffer_1608 = _RAND_1615[7:0];
  _RAND_1616 = {1{`RANDOM}};
  lineBuffer_1609 = _RAND_1616[7:0];
  _RAND_1617 = {1{`RANDOM}};
  lineBuffer_1610 = _RAND_1617[7:0];
  _RAND_1618 = {1{`RANDOM}};
  lineBuffer_1611 = _RAND_1618[7:0];
  _RAND_1619 = {1{`RANDOM}};
  lineBuffer_1612 = _RAND_1619[7:0];
  _RAND_1620 = {1{`RANDOM}};
  lineBuffer_1613 = _RAND_1620[7:0];
  _RAND_1621 = {1{`RANDOM}};
  lineBuffer_1614 = _RAND_1621[7:0];
  _RAND_1622 = {1{`RANDOM}};
  lineBuffer_1615 = _RAND_1622[7:0];
  _RAND_1623 = {1{`RANDOM}};
  lineBuffer_1616 = _RAND_1623[7:0];
  _RAND_1624 = {1{`RANDOM}};
  lineBuffer_1617 = _RAND_1624[7:0];
  _RAND_1625 = {1{`RANDOM}};
  lineBuffer_1618 = _RAND_1625[7:0];
  _RAND_1626 = {1{`RANDOM}};
  lineBuffer_1619 = _RAND_1626[7:0];
  _RAND_1627 = {1{`RANDOM}};
  lineBuffer_1620 = _RAND_1627[7:0];
  _RAND_1628 = {1{`RANDOM}};
  lineBuffer_1621 = _RAND_1628[7:0];
  _RAND_1629 = {1{`RANDOM}};
  lineBuffer_1622 = _RAND_1629[7:0];
  _RAND_1630 = {1{`RANDOM}};
  lineBuffer_1623 = _RAND_1630[7:0];
  _RAND_1631 = {1{`RANDOM}};
  lineBuffer_1624 = _RAND_1631[7:0];
  _RAND_1632 = {1{`RANDOM}};
  lineBuffer_1625 = _RAND_1632[7:0];
  _RAND_1633 = {1{`RANDOM}};
  lineBuffer_1626 = _RAND_1633[7:0];
  _RAND_1634 = {1{`RANDOM}};
  lineBuffer_1627 = _RAND_1634[7:0];
  _RAND_1635 = {1{`RANDOM}};
  lineBuffer_1628 = _RAND_1635[7:0];
  _RAND_1636 = {1{`RANDOM}};
  lineBuffer_1629 = _RAND_1636[7:0];
  _RAND_1637 = {1{`RANDOM}};
  lineBuffer_1630 = _RAND_1637[7:0];
  _RAND_1638 = {1{`RANDOM}};
  lineBuffer_1631 = _RAND_1638[7:0];
  _RAND_1639 = {1{`RANDOM}};
  lineBuffer_1632 = _RAND_1639[7:0];
  _RAND_1640 = {1{`RANDOM}};
  lineBuffer_1633 = _RAND_1640[7:0];
  _RAND_1641 = {1{`RANDOM}};
  lineBuffer_1634 = _RAND_1641[7:0];
  _RAND_1642 = {1{`RANDOM}};
  lineBuffer_1635 = _RAND_1642[7:0];
  _RAND_1643 = {1{`RANDOM}};
  lineBuffer_1636 = _RAND_1643[7:0];
  _RAND_1644 = {1{`RANDOM}};
  lineBuffer_1637 = _RAND_1644[7:0];
  _RAND_1645 = {1{`RANDOM}};
  lineBuffer_1638 = _RAND_1645[7:0];
  _RAND_1646 = {1{`RANDOM}};
  lineBuffer_1639 = _RAND_1646[7:0];
  _RAND_1647 = {1{`RANDOM}};
  lineBuffer_1640 = _RAND_1647[7:0];
  _RAND_1648 = {1{`RANDOM}};
  lineBuffer_1641 = _RAND_1648[7:0];
  _RAND_1649 = {1{`RANDOM}};
  lineBuffer_1642 = _RAND_1649[7:0];
  _RAND_1650 = {1{`RANDOM}};
  lineBuffer_1643 = _RAND_1650[7:0];
  _RAND_1651 = {1{`RANDOM}};
  lineBuffer_1644 = _RAND_1651[7:0];
  _RAND_1652 = {1{`RANDOM}};
  lineBuffer_1645 = _RAND_1652[7:0];
  _RAND_1653 = {1{`RANDOM}};
  lineBuffer_1646 = _RAND_1653[7:0];
  _RAND_1654 = {1{`RANDOM}};
  lineBuffer_1647 = _RAND_1654[7:0];
  _RAND_1655 = {1{`RANDOM}};
  lineBuffer_1648 = _RAND_1655[7:0];
  _RAND_1656 = {1{`RANDOM}};
  lineBuffer_1649 = _RAND_1656[7:0];
  _RAND_1657 = {1{`RANDOM}};
  lineBuffer_1650 = _RAND_1657[7:0];
  _RAND_1658 = {1{`RANDOM}};
  lineBuffer_1651 = _RAND_1658[7:0];
  _RAND_1659 = {1{`RANDOM}};
  lineBuffer_1652 = _RAND_1659[7:0];
  _RAND_1660 = {1{`RANDOM}};
  lineBuffer_1653 = _RAND_1660[7:0];
  _RAND_1661 = {1{`RANDOM}};
  lineBuffer_1654 = _RAND_1661[7:0];
  _RAND_1662 = {1{`RANDOM}};
  lineBuffer_1655 = _RAND_1662[7:0];
  _RAND_1663 = {1{`RANDOM}};
  lineBuffer_1656 = _RAND_1663[7:0];
  _RAND_1664 = {1{`RANDOM}};
  lineBuffer_1657 = _RAND_1664[7:0];
  _RAND_1665 = {1{`RANDOM}};
  lineBuffer_1658 = _RAND_1665[7:0];
  _RAND_1666 = {1{`RANDOM}};
  lineBuffer_1659 = _RAND_1666[7:0];
  _RAND_1667 = {1{`RANDOM}};
  lineBuffer_1660 = _RAND_1667[7:0];
  _RAND_1668 = {1{`RANDOM}};
  lineBuffer_1661 = _RAND_1668[7:0];
  _RAND_1669 = {1{`RANDOM}};
  lineBuffer_1662 = _RAND_1669[7:0];
  _RAND_1670 = {1{`RANDOM}};
  lineBuffer_1663 = _RAND_1670[7:0];
  _RAND_1671 = {1{`RANDOM}};
  lineBuffer_1664 = _RAND_1671[7:0];
  _RAND_1672 = {1{`RANDOM}};
  lineBuffer_1665 = _RAND_1672[7:0];
  _RAND_1673 = {1{`RANDOM}};
  lineBuffer_1666 = _RAND_1673[7:0];
  _RAND_1674 = {1{`RANDOM}};
  lineBuffer_1667 = _RAND_1674[7:0];
  _RAND_1675 = {1{`RANDOM}};
  lineBuffer_1668 = _RAND_1675[7:0];
  _RAND_1676 = {1{`RANDOM}};
  lineBuffer_1669 = _RAND_1676[7:0];
  _RAND_1677 = {1{`RANDOM}};
  lineBuffer_1670 = _RAND_1677[7:0];
  _RAND_1678 = {1{`RANDOM}};
  lineBuffer_1671 = _RAND_1678[7:0];
  _RAND_1679 = {1{`RANDOM}};
  lineBuffer_1672 = _RAND_1679[7:0];
  _RAND_1680 = {1{`RANDOM}};
  lineBuffer_1673 = _RAND_1680[7:0];
  _RAND_1681 = {1{`RANDOM}};
  lineBuffer_1674 = _RAND_1681[7:0];
  _RAND_1682 = {1{`RANDOM}};
  lineBuffer_1675 = _RAND_1682[7:0];
  _RAND_1683 = {1{`RANDOM}};
  lineBuffer_1676 = _RAND_1683[7:0];
  _RAND_1684 = {1{`RANDOM}};
  lineBuffer_1677 = _RAND_1684[7:0];
  _RAND_1685 = {1{`RANDOM}};
  lineBuffer_1678 = _RAND_1685[7:0];
  _RAND_1686 = {1{`RANDOM}};
  lineBuffer_1679 = _RAND_1686[7:0];
  _RAND_1687 = {1{`RANDOM}};
  lineBuffer_1680 = _RAND_1687[7:0];
  _RAND_1688 = {1{`RANDOM}};
  lineBuffer_1681 = _RAND_1688[7:0];
  _RAND_1689 = {1{`RANDOM}};
  lineBuffer_1682 = _RAND_1689[7:0];
  _RAND_1690 = {1{`RANDOM}};
  lineBuffer_1683 = _RAND_1690[7:0];
  _RAND_1691 = {1{`RANDOM}};
  lineBuffer_1684 = _RAND_1691[7:0];
  _RAND_1692 = {1{`RANDOM}};
  lineBuffer_1685 = _RAND_1692[7:0];
  _RAND_1693 = {1{`RANDOM}};
  lineBuffer_1686 = _RAND_1693[7:0];
  _RAND_1694 = {1{`RANDOM}};
  lineBuffer_1687 = _RAND_1694[7:0];
  _RAND_1695 = {1{`RANDOM}};
  lineBuffer_1688 = _RAND_1695[7:0];
  _RAND_1696 = {1{`RANDOM}};
  lineBuffer_1689 = _RAND_1696[7:0];
  _RAND_1697 = {1{`RANDOM}};
  lineBuffer_1690 = _RAND_1697[7:0];
  _RAND_1698 = {1{`RANDOM}};
  lineBuffer_1691 = _RAND_1698[7:0];
  _RAND_1699 = {1{`RANDOM}};
  lineBuffer_1692 = _RAND_1699[7:0];
  _RAND_1700 = {1{`RANDOM}};
  lineBuffer_1693 = _RAND_1700[7:0];
  _RAND_1701 = {1{`RANDOM}};
  lineBuffer_1694 = _RAND_1701[7:0];
  _RAND_1702 = {1{`RANDOM}};
  lineBuffer_1695 = _RAND_1702[7:0];
  _RAND_1703 = {1{`RANDOM}};
  lineBuffer_1696 = _RAND_1703[7:0];
  _RAND_1704 = {1{`RANDOM}};
  lineBuffer_1697 = _RAND_1704[7:0];
  _RAND_1705 = {1{`RANDOM}};
  lineBuffer_1698 = _RAND_1705[7:0];
  _RAND_1706 = {1{`RANDOM}};
  lineBuffer_1699 = _RAND_1706[7:0];
  _RAND_1707 = {1{`RANDOM}};
  lineBuffer_1700 = _RAND_1707[7:0];
  _RAND_1708 = {1{`RANDOM}};
  lineBuffer_1701 = _RAND_1708[7:0];
  _RAND_1709 = {1{`RANDOM}};
  lineBuffer_1702 = _RAND_1709[7:0];
  _RAND_1710 = {1{`RANDOM}};
  lineBuffer_1703 = _RAND_1710[7:0];
  _RAND_1711 = {1{`RANDOM}};
  lineBuffer_1704 = _RAND_1711[7:0];
  _RAND_1712 = {1{`RANDOM}};
  lineBuffer_1705 = _RAND_1712[7:0];
  _RAND_1713 = {1{`RANDOM}};
  lineBuffer_1706 = _RAND_1713[7:0];
  _RAND_1714 = {1{`RANDOM}};
  lineBuffer_1707 = _RAND_1714[7:0];
  _RAND_1715 = {1{`RANDOM}};
  lineBuffer_1708 = _RAND_1715[7:0];
  _RAND_1716 = {1{`RANDOM}};
  lineBuffer_1709 = _RAND_1716[7:0];
  _RAND_1717 = {1{`RANDOM}};
  lineBuffer_1710 = _RAND_1717[7:0];
  _RAND_1718 = {1{`RANDOM}};
  lineBuffer_1711 = _RAND_1718[7:0];
  _RAND_1719 = {1{`RANDOM}};
  lineBuffer_1712 = _RAND_1719[7:0];
  _RAND_1720 = {1{`RANDOM}};
  lineBuffer_1713 = _RAND_1720[7:0];
  _RAND_1721 = {1{`RANDOM}};
  lineBuffer_1714 = _RAND_1721[7:0];
  _RAND_1722 = {1{`RANDOM}};
  lineBuffer_1715 = _RAND_1722[7:0];
  _RAND_1723 = {1{`RANDOM}};
  lineBuffer_1716 = _RAND_1723[7:0];
  _RAND_1724 = {1{`RANDOM}};
  lineBuffer_1717 = _RAND_1724[7:0];
  _RAND_1725 = {1{`RANDOM}};
  lineBuffer_1718 = _RAND_1725[7:0];
  _RAND_1726 = {1{`RANDOM}};
  lineBuffer_1719 = _RAND_1726[7:0];
  _RAND_1727 = {1{`RANDOM}};
  lineBuffer_1720 = _RAND_1727[7:0];
  _RAND_1728 = {1{`RANDOM}};
  lineBuffer_1721 = _RAND_1728[7:0];
  _RAND_1729 = {1{`RANDOM}};
  lineBuffer_1722 = _RAND_1729[7:0];
  _RAND_1730 = {1{`RANDOM}};
  lineBuffer_1723 = _RAND_1730[7:0];
  _RAND_1731 = {1{`RANDOM}};
  lineBuffer_1724 = _RAND_1731[7:0];
  _RAND_1732 = {1{`RANDOM}};
  lineBuffer_1725 = _RAND_1732[7:0];
  _RAND_1733 = {1{`RANDOM}};
  lineBuffer_1726 = _RAND_1733[7:0];
  _RAND_1734 = {1{`RANDOM}};
  lineBuffer_1727 = _RAND_1734[7:0];
  _RAND_1735 = {1{`RANDOM}};
  lineBuffer_1728 = _RAND_1735[7:0];
  _RAND_1736 = {1{`RANDOM}};
  lineBuffer_1729 = _RAND_1736[7:0];
  _RAND_1737 = {1{`RANDOM}};
  lineBuffer_1730 = _RAND_1737[7:0];
  _RAND_1738 = {1{`RANDOM}};
  lineBuffer_1731 = _RAND_1738[7:0];
  _RAND_1739 = {1{`RANDOM}};
  lineBuffer_1732 = _RAND_1739[7:0];
  _RAND_1740 = {1{`RANDOM}};
  lineBuffer_1733 = _RAND_1740[7:0];
  _RAND_1741 = {1{`RANDOM}};
  lineBuffer_1734 = _RAND_1741[7:0];
  _RAND_1742 = {1{`RANDOM}};
  lineBuffer_1735 = _RAND_1742[7:0];
  _RAND_1743 = {1{`RANDOM}};
  lineBuffer_1736 = _RAND_1743[7:0];
  _RAND_1744 = {1{`RANDOM}};
  lineBuffer_1737 = _RAND_1744[7:0];
  _RAND_1745 = {1{`RANDOM}};
  lineBuffer_1738 = _RAND_1745[7:0];
  _RAND_1746 = {1{`RANDOM}};
  lineBuffer_1739 = _RAND_1746[7:0];
  _RAND_1747 = {1{`RANDOM}};
  lineBuffer_1740 = _RAND_1747[7:0];
  _RAND_1748 = {1{`RANDOM}};
  lineBuffer_1741 = _RAND_1748[7:0];
  _RAND_1749 = {1{`RANDOM}};
  lineBuffer_1742 = _RAND_1749[7:0];
  _RAND_1750 = {1{`RANDOM}};
  lineBuffer_1743 = _RAND_1750[7:0];
  _RAND_1751 = {1{`RANDOM}};
  lineBuffer_1744 = _RAND_1751[7:0];
  _RAND_1752 = {1{`RANDOM}};
  lineBuffer_1745 = _RAND_1752[7:0];
  _RAND_1753 = {1{`RANDOM}};
  lineBuffer_1746 = _RAND_1753[7:0];
  _RAND_1754 = {1{`RANDOM}};
  lineBuffer_1747 = _RAND_1754[7:0];
  _RAND_1755 = {1{`RANDOM}};
  lineBuffer_1748 = _RAND_1755[7:0];
  _RAND_1756 = {1{`RANDOM}};
  lineBuffer_1749 = _RAND_1756[7:0];
  _RAND_1757 = {1{`RANDOM}};
  lineBuffer_1750 = _RAND_1757[7:0];
  _RAND_1758 = {1{`RANDOM}};
  lineBuffer_1751 = _RAND_1758[7:0];
  _RAND_1759 = {1{`RANDOM}};
  lineBuffer_1752 = _RAND_1759[7:0];
  _RAND_1760 = {1{`RANDOM}};
  lineBuffer_1753 = _RAND_1760[7:0];
  _RAND_1761 = {1{`RANDOM}};
  lineBuffer_1754 = _RAND_1761[7:0];
  _RAND_1762 = {1{`RANDOM}};
  lineBuffer_1755 = _RAND_1762[7:0];
  _RAND_1763 = {1{`RANDOM}};
  lineBuffer_1756 = _RAND_1763[7:0];
  _RAND_1764 = {1{`RANDOM}};
  lineBuffer_1757 = _RAND_1764[7:0];
  _RAND_1765 = {1{`RANDOM}};
  lineBuffer_1758 = _RAND_1765[7:0];
  _RAND_1766 = {1{`RANDOM}};
  lineBuffer_1759 = _RAND_1766[7:0];
  _RAND_1767 = {1{`RANDOM}};
  lineBuffer_1760 = _RAND_1767[7:0];
  _RAND_1768 = {1{`RANDOM}};
  lineBuffer_1761 = _RAND_1768[7:0];
  _RAND_1769 = {1{`RANDOM}};
  lineBuffer_1762 = _RAND_1769[7:0];
  _RAND_1770 = {1{`RANDOM}};
  lineBuffer_1763 = _RAND_1770[7:0];
  _RAND_1771 = {1{`RANDOM}};
  lineBuffer_1764 = _RAND_1771[7:0];
  _RAND_1772 = {1{`RANDOM}};
  lineBuffer_1765 = _RAND_1772[7:0];
  _RAND_1773 = {1{`RANDOM}};
  lineBuffer_1766 = _RAND_1773[7:0];
  _RAND_1774 = {1{`RANDOM}};
  lineBuffer_1767 = _RAND_1774[7:0];
  _RAND_1775 = {1{`RANDOM}};
  lineBuffer_1768 = _RAND_1775[7:0];
  _RAND_1776 = {1{`RANDOM}};
  lineBuffer_1769 = _RAND_1776[7:0];
  _RAND_1777 = {1{`RANDOM}};
  lineBuffer_1770 = _RAND_1777[7:0];
  _RAND_1778 = {1{`RANDOM}};
  lineBuffer_1771 = _RAND_1778[7:0];
  _RAND_1779 = {1{`RANDOM}};
  lineBuffer_1772 = _RAND_1779[7:0];
  _RAND_1780 = {1{`RANDOM}};
  lineBuffer_1773 = _RAND_1780[7:0];
  _RAND_1781 = {1{`RANDOM}};
  lineBuffer_1774 = _RAND_1781[7:0];
  _RAND_1782 = {1{`RANDOM}};
  lineBuffer_1775 = _RAND_1782[7:0];
  _RAND_1783 = {1{`RANDOM}};
  lineBuffer_1776 = _RAND_1783[7:0];
  _RAND_1784 = {1{`RANDOM}};
  lineBuffer_1777 = _RAND_1784[7:0];
  _RAND_1785 = {1{`RANDOM}};
  lineBuffer_1778 = _RAND_1785[7:0];
  _RAND_1786 = {1{`RANDOM}};
  lineBuffer_1779 = _RAND_1786[7:0];
  _RAND_1787 = {1{`RANDOM}};
  lineBuffer_1780 = _RAND_1787[7:0];
  _RAND_1788 = {1{`RANDOM}};
  lineBuffer_1781 = _RAND_1788[7:0];
  _RAND_1789 = {1{`RANDOM}};
  lineBuffer_1782 = _RAND_1789[7:0];
  _RAND_1790 = {1{`RANDOM}};
  lineBuffer_1783 = _RAND_1790[7:0];
  _RAND_1791 = {1{`RANDOM}};
  lineBuffer_1784 = _RAND_1791[7:0];
  _RAND_1792 = {1{`RANDOM}};
  lineBuffer_1785 = _RAND_1792[7:0];
  _RAND_1793 = {1{`RANDOM}};
  lineBuffer_1786 = _RAND_1793[7:0];
  _RAND_1794 = {1{`RANDOM}};
  lineBuffer_1787 = _RAND_1794[7:0];
  _RAND_1795 = {1{`RANDOM}};
  lineBuffer_1788 = _RAND_1795[7:0];
  _RAND_1796 = {1{`RANDOM}};
  lineBuffer_1789 = _RAND_1796[7:0];
  _RAND_1797 = {1{`RANDOM}};
  lineBuffer_1790 = _RAND_1797[7:0];
  _RAND_1798 = {1{`RANDOM}};
  lineBuffer_1791 = _RAND_1798[7:0];
  _RAND_1799 = {1{`RANDOM}};
  lineBuffer_1792 = _RAND_1799[7:0];
  _RAND_1800 = {1{`RANDOM}};
  lineBuffer_1793 = _RAND_1800[7:0];
  _RAND_1801 = {1{`RANDOM}};
  lineBuffer_1794 = _RAND_1801[7:0];
  _RAND_1802 = {1{`RANDOM}};
  lineBuffer_1795 = _RAND_1802[7:0];
  _RAND_1803 = {1{`RANDOM}};
  lineBuffer_1796 = _RAND_1803[7:0];
  _RAND_1804 = {1{`RANDOM}};
  lineBuffer_1797 = _RAND_1804[7:0];
  _RAND_1805 = {1{`RANDOM}};
  lineBuffer_1798 = _RAND_1805[7:0];
  _RAND_1806 = {1{`RANDOM}};
  lineBuffer_1799 = _RAND_1806[7:0];
  _RAND_1807 = {1{`RANDOM}};
  lineBuffer_1800 = _RAND_1807[7:0];
  _RAND_1808 = {1{`RANDOM}};
  lineBuffer_1801 = _RAND_1808[7:0];
  _RAND_1809 = {1{`RANDOM}};
  lineBuffer_1802 = _RAND_1809[7:0];
  _RAND_1810 = {1{`RANDOM}};
  lineBuffer_1803 = _RAND_1810[7:0];
  _RAND_1811 = {1{`RANDOM}};
  lineBuffer_1804 = _RAND_1811[7:0];
  _RAND_1812 = {1{`RANDOM}};
  lineBuffer_1805 = _RAND_1812[7:0];
  _RAND_1813 = {1{`RANDOM}};
  lineBuffer_1806 = _RAND_1813[7:0];
  _RAND_1814 = {1{`RANDOM}};
  lineBuffer_1807 = _RAND_1814[7:0];
  _RAND_1815 = {1{`RANDOM}};
  lineBuffer_1808 = _RAND_1815[7:0];
  _RAND_1816 = {1{`RANDOM}};
  lineBuffer_1809 = _RAND_1816[7:0];
  _RAND_1817 = {1{`RANDOM}};
  lineBuffer_1810 = _RAND_1817[7:0];
  _RAND_1818 = {1{`RANDOM}};
  lineBuffer_1811 = _RAND_1818[7:0];
  _RAND_1819 = {1{`RANDOM}};
  lineBuffer_1812 = _RAND_1819[7:0];
  _RAND_1820 = {1{`RANDOM}};
  lineBuffer_1813 = _RAND_1820[7:0];
  _RAND_1821 = {1{`RANDOM}};
  lineBuffer_1814 = _RAND_1821[7:0];
  _RAND_1822 = {1{`RANDOM}};
  lineBuffer_1815 = _RAND_1822[7:0];
  _RAND_1823 = {1{`RANDOM}};
  lineBuffer_1816 = _RAND_1823[7:0];
  _RAND_1824 = {1{`RANDOM}};
  lineBuffer_1817 = _RAND_1824[7:0];
  _RAND_1825 = {1{`RANDOM}};
  lineBuffer_1818 = _RAND_1825[7:0];
  _RAND_1826 = {1{`RANDOM}};
  lineBuffer_1819 = _RAND_1826[7:0];
  _RAND_1827 = {1{`RANDOM}};
  lineBuffer_1820 = _RAND_1827[7:0];
  _RAND_1828 = {1{`RANDOM}};
  lineBuffer_1821 = _RAND_1828[7:0];
  _RAND_1829 = {1{`RANDOM}};
  lineBuffer_1822 = _RAND_1829[7:0];
  _RAND_1830 = {1{`RANDOM}};
  lineBuffer_1823 = _RAND_1830[7:0];
  _RAND_1831 = {1{`RANDOM}};
  lineBuffer_1824 = _RAND_1831[7:0];
  _RAND_1832 = {1{`RANDOM}};
  lineBuffer_1825 = _RAND_1832[7:0];
  _RAND_1833 = {1{`RANDOM}};
  lineBuffer_1826 = _RAND_1833[7:0];
  _RAND_1834 = {1{`RANDOM}};
  lineBuffer_1827 = _RAND_1834[7:0];
  _RAND_1835 = {1{`RANDOM}};
  lineBuffer_1828 = _RAND_1835[7:0];
  _RAND_1836 = {1{`RANDOM}};
  lineBuffer_1829 = _RAND_1836[7:0];
  _RAND_1837 = {1{`RANDOM}};
  lineBuffer_1830 = _RAND_1837[7:0];
  _RAND_1838 = {1{`RANDOM}};
  lineBuffer_1831 = _RAND_1838[7:0];
  _RAND_1839 = {1{`RANDOM}};
  lineBuffer_1832 = _RAND_1839[7:0];
  _RAND_1840 = {1{`RANDOM}};
  lineBuffer_1833 = _RAND_1840[7:0];
  _RAND_1841 = {1{`RANDOM}};
  lineBuffer_1834 = _RAND_1841[7:0];
  _RAND_1842 = {1{`RANDOM}};
  lineBuffer_1835 = _RAND_1842[7:0];
  _RAND_1843 = {1{`RANDOM}};
  lineBuffer_1836 = _RAND_1843[7:0];
  _RAND_1844 = {1{`RANDOM}};
  lineBuffer_1837 = _RAND_1844[7:0];
  _RAND_1845 = {1{`RANDOM}};
  lineBuffer_1838 = _RAND_1845[7:0];
  _RAND_1846 = {1{`RANDOM}};
  lineBuffer_1839 = _RAND_1846[7:0];
  _RAND_1847 = {1{`RANDOM}};
  lineBuffer_1840 = _RAND_1847[7:0];
  _RAND_1848 = {1{`RANDOM}};
  lineBuffer_1841 = _RAND_1848[7:0];
  _RAND_1849 = {1{`RANDOM}};
  lineBuffer_1842 = _RAND_1849[7:0];
  _RAND_1850 = {1{`RANDOM}};
  lineBuffer_1843 = _RAND_1850[7:0];
  _RAND_1851 = {1{`RANDOM}};
  lineBuffer_1844 = _RAND_1851[7:0];
  _RAND_1852 = {1{`RANDOM}};
  lineBuffer_1845 = _RAND_1852[7:0];
  _RAND_1853 = {1{`RANDOM}};
  lineBuffer_1846 = _RAND_1853[7:0];
  _RAND_1854 = {1{`RANDOM}};
  lineBuffer_1847 = _RAND_1854[7:0];
  _RAND_1855 = {1{`RANDOM}};
  lineBuffer_1848 = _RAND_1855[7:0];
  _RAND_1856 = {1{`RANDOM}};
  lineBuffer_1849 = _RAND_1856[7:0];
  _RAND_1857 = {1{`RANDOM}};
  lineBuffer_1850 = _RAND_1857[7:0];
  _RAND_1858 = {1{`RANDOM}};
  lineBuffer_1851 = _RAND_1858[7:0];
  _RAND_1859 = {1{`RANDOM}};
  lineBuffer_1852 = _RAND_1859[7:0];
  _RAND_1860 = {1{`RANDOM}};
  lineBuffer_1853 = _RAND_1860[7:0];
  _RAND_1861 = {1{`RANDOM}};
  lineBuffer_1854 = _RAND_1861[7:0];
  _RAND_1862 = {1{`RANDOM}};
  lineBuffer_1855 = _RAND_1862[7:0];
  _RAND_1863 = {1{`RANDOM}};
  lineBuffer_1856 = _RAND_1863[7:0];
  _RAND_1864 = {1{`RANDOM}};
  lineBuffer_1857 = _RAND_1864[7:0];
  _RAND_1865 = {1{`RANDOM}};
  lineBuffer_1858 = _RAND_1865[7:0];
  _RAND_1866 = {1{`RANDOM}};
  lineBuffer_1859 = _RAND_1866[7:0];
  _RAND_1867 = {1{`RANDOM}};
  lineBuffer_1860 = _RAND_1867[7:0];
  _RAND_1868 = {1{`RANDOM}};
  lineBuffer_1861 = _RAND_1868[7:0];
  _RAND_1869 = {1{`RANDOM}};
  lineBuffer_1862 = _RAND_1869[7:0];
  _RAND_1870 = {1{`RANDOM}};
  lineBuffer_1863 = _RAND_1870[7:0];
  _RAND_1871 = {1{`RANDOM}};
  lineBuffer_1864 = _RAND_1871[7:0];
  _RAND_1872 = {1{`RANDOM}};
  lineBuffer_1865 = _RAND_1872[7:0];
  _RAND_1873 = {1{`RANDOM}};
  lineBuffer_1866 = _RAND_1873[7:0];
  _RAND_1874 = {1{`RANDOM}};
  lineBuffer_1867 = _RAND_1874[7:0];
  _RAND_1875 = {1{`RANDOM}};
  lineBuffer_1868 = _RAND_1875[7:0];
  _RAND_1876 = {1{`RANDOM}};
  lineBuffer_1869 = _RAND_1876[7:0];
  _RAND_1877 = {1{`RANDOM}};
  lineBuffer_1870 = _RAND_1877[7:0];
  _RAND_1878 = {1{`RANDOM}};
  lineBuffer_1871 = _RAND_1878[7:0];
  _RAND_1879 = {1{`RANDOM}};
  lineBuffer_1872 = _RAND_1879[7:0];
  _RAND_1880 = {1{`RANDOM}};
  lineBuffer_1873 = _RAND_1880[7:0];
  _RAND_1881 = {1{`RANDOM}};
  lineBuffer_1874 = _RAND_1881[7:0];
  _RAND_1882 = {1{`RANDOM}};
  lineBuffer_1875 = _RAND_1882[7:0];
  _RAND_1883 = {1{`RANDOM}};
  lineBuffer_1876 = _RAND_1883[7:0];
  _RAND_1884 = {1{`RANDOM}};
  lineBuffer_1877 = _RAND_1884[7:0];
  _RAND_1885 = {1{`RANDOM}};
  lineBuffer_1878 = _RAND_1885[7:0];
  _RAND_1886 = {1{`RANDOM}};
  lineBuffer_1879 = _RAND_1886[7:0];
  _RAND_1887 = {1{`RANDOM}};
  lineBuffer_1880 = _RAND_1887[7:0];
  _RAND_1888 = {1{`RANDOM}};
  lineBuffer_1881 = _RAND_1888[7:0];
  _RAND_1889 = {1{`RANDOM}};
  lineBuffer_1882 = _RAND_1889[7:0];
  _RAND_1890 = {1{`RANDOM}};
  lineBuffer_1883 = _RAND_1890[7:0];
  _RAND_1891 = {1{`RANDOM}};
  lineBuffer_1884 = _RAND_1891[7:0];
  _RAND_1892 = {1{`RANDOM}};
  lineBuffer_1885 = _RAND_1892[7:0];
  _RAND_1893 = {1{`RANDOM}};
  lineBuffer_1886 = _RAND_1893[7:0];
  _RAND_1894 = {1{`RANDOM}};
  lineBuffer_1887 = _RAND_1894[7:0];
  _RAND_1895 = {1{`RANDOM}};
  lineBuffer_1888 = _RAND_1895[7:0];
  _RAND_1896 = {1{`RANDOM}};
  lineBuffer_1889 = _RAND_1896[7:0];
  _RAND_1897 = {1{`RANDOM}};
  lineBuffer_1890 = _RAND_1897[7:0];
  _RAND_1898 = {1{`RANDOM}};
  lineBuffer_1891 = _RAND_1898[7:0];
  _RAND_1899 = {1{`RANDOM}};
  lineBuffer_1892 = _RAND_1899[7:0];
  _RAND_1900 = {1{`RANDOM}};
  lineBuffer_1893 = _RAND_1900[7:0];
  _RAND_1901 = {1{`RANDOM}};
  lineBuffer_1894 = _RAND_1901[7:0];
  _RAND_1902 = {1{`RANDOM}};
  lineBuffer_1895 = _RAND_1902[7:0];
  _RAND_1903 = {1{`RANDOM}};
  lineBuffer_1896 = _RAND_1903[7:0];
  _RAND_1904 = {1{`RANDOM}};
  lineBuffer_1897 = _RAND_1904[7:0];
  _RAND_1905 = {1{`RANDOM}};
  lineBuffer_1898 = _RAND_1905[7:0];
  _RAND_1906 = {1{`RANDOM}};
  lineBuffer_1899 = _RAND_1906[7:0];
  _RAND_1907 = {1{`RANDOM}};
  lineBuffer_1900 = _RAND_1907[7:0];
  _RAND_1908 = {1{`RANDOM}};
  lineBuffer_1901 = _RAND_1908[7:0];
  _RAND_1909 = {1{`RANDOM}};
  lineBuffer_1902 = _RAND_1909[7:0];
  _RAND_1910 = {1{`RANDOM}};
  lineBuffer_1903 = _RAND_1910[7:0];
  _RAND_1911 = {1{`RANDOM}};
  lineBuffer_1904 = _RAND_1911[7:0];
  _RAND_1912 = {1{`RANDOM}};
  lineBuffer_1905 = _RAND_1912[7:0];
  _RAND_1913 = {1{`RANDOM}};
  lineBuffer_1906 = _RAND_1913[7:0];
  _RAND_1914 = {1{`RANDOM}};
  lineBuffer_1907 = _RAND_1914[7:0];
  _RAND_1915 = {1{`RANDOM}};
  lineBuffer_1908 = _RAND_1915[7:0];
  _RAND_1916 = {1{`RANDOM}};
  lineBuffer_1909 = _RAND_1916[7:0];
  _RAND_1917 = {1{`RANDOM}};
  lineBuffer_1910 = _RAND_1917[7:0];
  _RAND_1918 = {1{`RANDOM}};
  lineBuffer_1911 = _RAND_1918[7:0];
  _RAND_1919 = {1{`RANDOM}};
  lineBuffer_1912 = _RAND_1919[7:0];
  _RAND_1920 = {1{`RANDOM}};
  lineBuffer_1913 = _RAND_1920[7:0];
  _RAND_1921 = {1{`RANDOM}};
  lineBuffer_1914 = _RAND_1921[7:0];
  _RAND_1922 = {1{`RANDOM}};
  lineBuffer_1915 = _RAND_1922[7:0];
  _RAND_1923 = {1{`RANDOM}};
  lineBuffer_1916 = _RAND_1923[7:0];
  _RAND_1924 = {1{`RANDOM}};
  lineBuffer_1917 = _RAND_1924[7:0];
  _RAND_1925 = {1{`RANDOM}};
  lineBuffer_1918 = _RAND_1925[7:0];
  _RAND_1926 = {1{`RANDOM}};
  lineBuffer_1919 = _RAND_1926[7:0];
  _RAND_1927 = {1{`RANDOM}};
  lineBuffer_1920 = _RAND_1927[7:0];
  _RAND_1928 = {1{`RANDOM}};
  lineBuffer_1921 = _RAND_1928[7:0];
  _RAND_1929 = {1{`RANDOM}};
  lineBuffer_1922 = _RAND_1929[7:0];
  _RAND_1930 = {1{`RANDOM}};
  lineBuffer_1923 = _RAND_1930[7:0];
  _RAND_1931 = {1{`RANDOM}};
  lineBuffer_1924 = _RAND_1931[7:0];
  _RAND_1932 = {1{`RANDOM}};
  lineBuffer_1925 = _RAND_1932[7:0];
  _RAND_1933 = {1{`RANDOM}};
  lineBuffer_1926 = _RAND_1933[7:0];
  _RAND_1934 = {1{`RANDOM}};
  lineBuffer_1927 = _RAND_1934[7:0];
  _RAND_1935 = {1{`RANDOM}};
  lineBuffer_1928 = _RAND_1935[7:0];
  _RAND_1936 = {1{`RANDOM}};
  lineBuffer_1929 = _RAND_1936[7:0];
  _RAND_1937 = {1{`RANDOM}};
  lineBuffer_1930 = _RAND_1937[7:0];
  _RAND_1938 = {1{`RANDOM}};
  lineBuffer_1931 = _RAND_1938[7:0];
  _RAND_1939 = {1{`RANDOM}};
  lineBuffer_1932 = _RAND_1939[7:0];
  _RAND_1940 = {1{`RANDOM}};
  lineBuffer_1933 = _RAND_1940[7:0];
  _RAND_1941 = {1{`RANDOM}};
  lineBuffer_1934 = _RAND_1941[7:0];
  _RAND_1942 = {1{`RANDOM}};
  lineBuffer_1935 = _RAND_1942[7:0];
  _RAND_1943 = {1{`RANDOM}};
  lineBuffer_1936 = _RAND_1943[7:0];
  _RAND_1944 = {1{`RANDOM}};
  lineBuffer_1937 = _RAND_1944[7:0];
  _RAND_1945 = {1{`RANDOM}};
  lineBuffer_1938 = _RAND_1945[7:0];
  _RAND_1946 = {1{`RANDOM}};
  lineBuffer_1939 = _RAND_1946[7:0];
  _RAND_1947 = {1{`RANDOM}};
  lineBuffer_1940 = _RAND_1947[7:0];
  _RAND_1948 = {1{`RANDOM}};
  lineBuffer_1941 = _RAND_1948[7:0];
  _RAND_1949 = {1{`RANDOM}};
  lineBuffer_1942 = _RAND_1949[7:0];
  _RAND_1950 = {1{`RANDOM}};
  lineBuffer_1943 = _RAND_1950[7:0];
  _RAND_1951 = {1{`RANDOM}};
  lineBuffer_1944 = _RAND_1951[7:0];
  _RAND_1952 = {1{`RANDOM}};
  lineBuffer_1945 = _RAND_1952[7:0];
  _RAND_1953 = {1{`RANDOM}};
  lineBuffer_1946 = _RAND_1953[7:0];
  _RAND_1954 = {1{`RANDOM}};
  lineBuffer_1947 = _RAND_1954[7:0];
  _RAND_1955 = {1{`RANDOM}};
  lineBuffer_1948 = _RAND_1955[7:0];
  _RAND_1956 = {1{`RANDOM}};
  lineBuffer_1949 = _RAND_1956[7:0];
  _RAND_1957 = {1{`RANDOM}};
  lineBuffer_1950 = _RAND_1957[7:0];
  _RAND_1958 = {1{`RANDOM}};
  lineBuffer_1951 = _RAND_1958[7:0];
  _RAND_1959 = {1{`RANDOM}};
  lineBuffer_1952 = _RAND_1959[7:0];
  _RAND_1960 = {1{`RANDOM}};
  lineBuffer_1953 = _RAND_1960[7:0];
  _RAND_1961 = {1{`RANDOM}};
  lineBuffer_1954 = _RAND_1961[7:0];
  _RAND_1962 = {1{`RANDOM}};
  lineBuffer_1955 = _RAND_1962[7:0];
  _RAND_1963 = {1{`RANDOM}};
  lineBuffer_1956 = _RAND_1963[7:0];
  _RAND_1964 = {1{`RANDOM}};
  lineBuffer_1957 = _RAND_1964[7:0];
  _RAND_1965 = {1{`RANDOM}};
  lineBuffer_1958 = _RAND_1965[7:0];
  _RAND_1966 = {1{`RANDOM}};
  lineBuffer_1959 = _RAND_1966[7:0];
  _RAND_1967 = {1{`RANDOM}};
  lineBuffer_1960 = _RAND_1967[7:0];
  _RAND_1968 = {1{`RANDOM}};
  lineBuffer_1961 = _RAND_1968[7:0];
  _RAND_1969 = {1{`RANDOM}};
  lineBuffer_1962 = _RAND_1969[7:0];
  _RAND_1970 = {1{`RANDOM}};
  lineBuffer_1963 = _RAND_1970[7:0];
  _RAND_1971 = {1{`RANDOM}};
  lineBuffer_1964 = _RAND_1971[7:0];
  _RAND_1972 = {1{`RANDOM}};
  lineBuffer_1965 = _RAND_1972[7:0];
  _RAND_1973 = {1{`RANDOM}};
  lineBuffer_1966 = _RAND_1973[7:0];
  _RAND_1974 = {1{`RANDOM}};
  lineBuffer_1967 = _RAND_1974[7:0];
  _RAND_1975 = {1{`RANDOM}};
  lineBuffer_1968 = _RAND_1975[7:0];
  _RAND_1976 = {1{`RANDOM}};
  lineBuffer_1969 = _RAND_1976[7:0];
  _RAND_1977 = {1{`RANDOM}};
  lineBuffer_1970 = _RAND_1977[7:0];
  _RAND_1978 = {1{`RANDOM}};
  lineBuffer_1971 = _RAND_1978[7:0];
  _RAND_1979 = {1{`RANDOM}};
  lineBuffer_1972 = _RAND_1979[7:0];
  _RAND_1980 = {1{`RANDOM}};
  lineBuffer_1973 = _RAND_1980[7:0];
  _RAND_1981 = {1{`RANDOM}};
  lineBuffer_1974 = _RAND_1981[7:0];
  _RAND_1982 = {1{`RANDOM}};
  lineBuffer_1975 = _RAND_1982[7:0];
  _RAND_1983 = {1{`RANDOM}};
  lineBuffer_1976 = _RAND_1983[7:0];
  _RAND_1984 = {1{`RANDOM}};
  lineBuffer_1977 = _RAND_1984[7:0];
  _RAND_1985 = {1{`RANDOM}};
  lineBuffer_1978 = _RAND_1985[7:0];
  _RAND_1986 = {1{`RANDOM}};
  lineBuffer_1979 = _RAND_1986[7:0];
  _RAND_1987 = {1{`RANDOM}};
  lineBuffer_1980 = _RAND_1987[7:0];
  _RAND_1988 = {1{`RANDOM}};
  lineBuffer_1981 = _RAND_1988[7:0];
  _RAND_1989 = {1{`RANDOM}};
  lineBuffer_1982 = _RAND_1989[7:0];
  _RAND_1990 = {1{`RANDOM}};
  lineBuffer_1983 = _RAND_1990[7:0];
  _RAND_1991 = {1{`RANDOM}};
  lineBuffer_1984 = _RAND_1991[7:0];
  _RAND_1992 = {1{`RANDOM}};
  lineBuffer_1985 = _RAND_1992[7:0];
  _RAND_1993 = {1{`RANDOM}};
  lineBuffer_1986 = _RAND_1993[7:0];
  _RAND_1994 = {1{`RANDOM}};
  lineBuffer_1987 = _RAND_1994[7:0];
  _RAND_1995 = {1{`RANDOM}};
  lineBuffer_1988 = _RAND_1995[7:0];
  _RAND_1996 = {1{`RANDOM}};
  lineBuffer_1989 = _RAND_1996[7:0];
  _RAND_1997 = {1{`RANDOM}};
  lineBuffer_1990 = _RAND_1997[7:0];
  _RAND_1998 = {1{`RANDOM}};
  lineBuffer_1991 = _RAND_1998[7:0];
  _RAND_1999 = {1{`RANDOM}};
  lineBuffer_1992 = _RAND_1999[7:0];
  _RAND_2000 = {1{`RANDOM}};
  lineBuffer_1993 = _RAND_2000[7:0];
  _RAND_2001 = {1{`RANDOM}};
  lineBuffer_1994 = _RAND_2001[7:0];
  _RAND_2002 = {1{`RANDOM}};
  lineBuffer_1995 = _RAND_2002[7:0];
  _RAND_2003 = {1{`RANDOM}};
  lineBuffer_1996 = _RAND_2003[7:0];
  _RAND_2004 = {1{`RANDOM}};
  lineBuffer_1997 = _RAND_2004[7:0];
  _RAND_2005 = {1{`RANDOM}};
  lineBuffer_1998 = _RAND_2005[7:0];
  _RAND_2006 = {1{`RANDOM}};
  lineBuffer_1999 = _RAND_2006[7:0];
  _RAND_2007 = {1{`RANDOM}};
  lineBuffer_2000 = _RAND_2007[7:0];
  _RAND_2008 = {1{`RANDOM}};
  lineBuffer_2001 = _RAND_2008[7:0];
  _RAND_2009 = {1{`RANDOM}};
  lineBuffer_2002 = _RAND_2009[7:0];
  _RAND_2010 = {1{`RANDOM}};
  lineBuffer_2003 = _RAND_2010[7:0];
  _RAND_2011 = {1{`RANDOM}};
  lineBuffer_2004 = _RAND_2011[7:0];
  _RAND_2012 = {1{`RANDOM}};
  lineBuffer_2005 = _RAND_2012[7:0];
  _RAND_2013 = {1{`RANDOM}};
  lineBuffer_2006 = _RAND_2013[7:0];
  _RAND_2014 = {1{`RANDOM}};
  lineBuffer_2007 = _RAND_2014[7:0];
  _RAND_2015 = {1{`RANDOM}};
  lineBuffer_2008 = _RAND_2015[7:0];
  _RAND_2016 = {1{`RANDOM}};
  lineBuffer_2009 = _RAND_2016[7:0];
  _RAND_2017 = {1{`RANDOM}};
  lineBuffer_2010 = _RAND_2017[7:0];
  _RAND_2018 = {1{`RANDOM}};
  lineBuffer_2011 = _RAND_2018[7:0];
  _RAND_2019 = {1{`RANDOM}};
  lineBuffer_2012 = _RAND_2019[7:0];
  _RAND_2020 = {1{`RANDOM}};
  lineBuffer_2013 = _RAND_2020[7:0];
  _RAND_2021 = {1{`RANDOM}};
  lineBuffer_2014 = _RAND_2021[7:0];
  _RAND_2022 = {1{`RANDOM}};
  lineBuffer_2015 = _RAND_2022[7:0];
  _RAND_2023 = {1{`RANDOM}};
  lineBuffer_2016 = _RAND_2023[7:0];
  _RAND_2024 = {1{`RANDOM}};
  lineBuffer_2017 = _RAND_2024[7:0];
  _RAND_2025 = {1{`RANDOM}};
  lineBuffer_2018 = _RAND_2025[7:0];
  _RAND_2026 = {1{`RANDOM}};
  lineBuffer_2019 = _RAND_2026[7:0];
  _RAND_2027 = {1{`RANDOM}};
  lineBuffer_2020 = _RAND_2027[7:0];
  _RAND_2028 = {1{`RANDOM}};
  lineBuffer_2021 = _RAND_2028[7:0];
  _RAND_2029 = {1{`RANDOM}};
  lineBuffer_2022 = _RAND_2029[7:0];
  _RAND_2030 = {1{`RANDOM}};
  lineBuffer_2023 = _RAND_2030[7:0];
  _RAND_2031 = {1{`RANDOM}};
  lineBuffer_2024 = _RAND_2031[7:0];
  _RAND_2032 = {1{`RANDOM}};
  lineBuffer_2025 = _RAND_2032[7:0];
  _RAND_2033 = {1{`RANDOM}};
  lineBuffer_2026 = _RAND_2033[7:0];
  _RAND_2034 = {1{`RANDOM}};
  lineBuffer_2027 = _RAND_2034[7:0];
  _RAND_2035 = {1{`RANDOM}};
  lineBuffer_2028 = _RAND_2035[7:0];
  _RAND_2036 = {1{`RANDOM}};
  lineBuffer_2029 = _RAND_2036[7:0];
  _RAND_2037 = {1{`RANDOM}};
  lineBuffer_2030 = _RAND_2037[7:0];
  _RAND_2038 = {1{`RANDOM}};
  lineBuffer_2031 = _RAND_2038[7:0];
  _RAND_2039 = {1{`RANDOM}};
  lineBuffer_2032 = _RAND_2039[7:0];
  _RAND_2040 = {1{`RANDOM}};
  lineBuffer_2033 = _RAND_2040[7:0];
  _RAND_2041 = {1{`RANDOM}};
  lineBuffer_2034 = _RAND_2041[7:0];
  _RAND_2042 = {1{`RANDOM}};
  lineBuffer_2035 = _RAND_2042[7:0];
  _RAND_2043 = {1{`RANDOM}};
  lineBuffer_2036 = _RAND_2043[7:0];
  _RAND_2044 = {1{`RANDOM}};
  lineBuffer_2037 = _RAND_2044[7:0];
  _RAND_2045 = {1{`RANDOM}};
  lineBuffer_2038 = _RAND_2045[7:0];
  _RAND_2046 = {1{`RANDOM}};
  lineBuffer_2039 = _RAND_2046[7:0];
  _RAND_2047 = {1{`RANDOM}};
  lineBuffer_2040 = _RAND_2047[7:0];
  _RAND_2048 = {1{`RANDOM}};
  lineBuffer_2041 = _RAND_2048[7:0];
  _RAND_2049 = {1{`RANDOM}};
  lineBuffer_2042 = _RAND_2049[7:0];
  _RAND_2050 = {1{`RANDOM}};
  lineBuffer_2043 = _RAND_2050[7:0];
  _RAND_2051 = {1{`RANDOM}};
  lineBuffer_2044 = _RAND_2051[7:0];
  _RAND_2052 = {1{`RANDOM}};
  lineBuffer_2045 = _RAND_2052[7:0];
  _RAND_2053 = {1{`RANDOM}};
  lineBuffer_2046 = _RAND_2053[7:0];
  _RAND_2054 = {1{`RANDOM}};
  lineBuffer_2047 = _RAND_2054[7:0];
  _RAND_2055 = {1{`RANDOM}};
  lineBuffer_2048 = _RAND_2055[7:0];
  _RAND_2056 = {1{`RANDOM}};
  lineBuffer_2049 = _RAND_2056[7:0];
  _RAND_2057 = {1{`RANDOM}};
  lineBuffer_2050 = _RAND_2057[7:0];
  _RAND_2058 = {1{`RANDOM}};
  lineBuffer_2051 = _RAND_2058[7:0];
  _RAND_2059 = {1{`RANDOM}};
  lineBuffer_2052 = _RAND_2059[7:0];
  _RAND_2060 = {1{`RANDOM}};
  lineBuffer_2053 = _RAND_2060[7:0];
  _RAND_2061 = {1{`RANDOM}};
  lineBuffer_2054 = _RAND_2061[7:0];
  _RAND_2062 = {1{`RANDOM}};
  lineBuffer_2055 = _RAND_2062[7:0];
  _RAND_2063 = {1{`RANDOM}};
  lineBuffer_2056 = _RAND_2063[7:0];
  _RAND_2064 = {1{`RANDOM}};
  lineBuffer_2057 = _RAND_2064[7:0];
  _RAND_2065 = {1{`RANDOM}};
  lineBuffer_2058 = _RAND_2065[7:0];
  _RAND_2066 = {1{`RANDOM}};
  lineBuffer_2059 = _RAND_2066[7:0];
  _RAND_2067 = {1{`RANDOM}};
  lineBuffer_2060 = _RAND_2067[7:0];
  _RAND_2068 = {1{`RANDOM}};
  lineBuffer_2061 = _RAND_2068[7:0];
  _RAND_2069 = {1{`RANDOM}};
  lineBuffer_2062 = _RAND_2069[7:0];
  _RAND_2070 = {1{`RANDOM}};
  lineBuffer_2063 = _RAND_2070[7:0];
  _RAND_2071 = {1{`RANDOM}};
  lineBuffer_2064 = _RAND_2071[7:0];
  _RAND_2072 = {1{`RANDOM}};
  lineBuffer_2065 = _RAND_2072[7:0];
  _RAND_2073 = {1{`RANDOM}};
  lineBuffer_2066 = _RAND_2073[7:0];
  _RAND_2074 = {1{`RANDOM}};
  lineBuffer_2067 = _RAND_2074[7:0];
  _RAND_2075 = {1{`RANDOM}};
  lineBuffer_2068 = _RAND_2075[7:0];
  _RAND_2076 = {1{`RANDOM}};
  lineBuffer_2069 = _RAND_2076[7:0];
  _RAND_2077 = {1{`RANDOM}};
  lineBuffer_2070 = _RAND_2077[7:0];
  _RAND_2078 = {1{`RANDOM}};
  lineBuffer_2071 = _RAND_2078[7:0];
  _RAND_2079 = {1{`RANDOM}};
  lineBuffer_2072 = _RAND_2079[7:0];
  _RAND_2080 = {1{`RANDOM}};
  lineBuffer_2073 = _RAND_2080[7:0];
  _RAND_2081 = {1{`RANDOM}};
  lineBuffer_2074 = _RAND_2081[7:0];
  _RAND_2082 = {1{`RANDOM}};
  lineBuffer_2075 = _RAND_2082[7:0];
  _RAND_2083 = {1{`RANDOM}};
  lineBuffer_2076 = _RAND_2083[7:0];
  _RAND_2084 = {1{`RANDOM}};
  lineBuffer_2077 = _RAND_2084[7:0];
  _RAND_2085 = {1{`RANDOM}};
  lineBuffer_2078 = _RAND_2085[7:0];
  _RAND_2086 = {1{`RANDOM}};
  lineBuffer_2079 = _RAND_2086[7:0];
  _RAND_2087 = {1{`RANDOM}};
  lineBuffer_2080 = _RAND_2087[7:0];
  _RAND_2088 = {1{`RANDOM}};
  lineBuffer_2081 = _RAND_2088[7:0];
  _RAND_2089 = {1{`RANDOM}};
  lineBuffer_2082 = _RAND_2089[7:0];
  _RAND_2090 = {1{`RANDOM}};
  lineBuffer_2083 = _RAND_2090[7:0];
  _RAND_2091 = {1{`RANDOM}};
  lineBuffer_2084 = _RAND_2091[7:0];
  _RAND_2092 = {1{`RANDOM}};
  lineBuffer_2085 = _RAND_2092[7:0];
  _RAND_2093 = {1{`RANDOM}};
  lineBuffer_2086 = _RAND_2093[7:0];
  _RAND_2094 = {1{`RANDOM}};
  lineBuffer_2087 = _RAND_2094[7:0];
  _RAND_2095 = {1{`RANDOM}};
  lineBuffer_2088 = _RAND_2095[7:0];
  _RAND_2096 = {1{`RANDOM}};
  lineBuffer_2089 = _RAND_2096[7:0];
  _RAND_2097 = {1{`RANDOM}};
  lineBuffer_2090 = _RAND_2097[7:0];
  _RAND_2098 = {1{`RANDOM}};
  lineBuffer_2091 = _RAND_2098[7:0];
  _RAND_2099 = {1{`RANDOM}};
  lineBuffer_2092 = _RAND_2099[7:0];
  _RAND_2100 = {1{`RANDOM}};
  lineBuffer_2093 = _RAND_2100[7:0];
  _RAND_2101 = {1{`RANDOM}};
  lineBuffer_2094 = _RAND_2101[7:0];
  _RAND_2102 = {1{`RANDOM}};
  lineBuffer_2095 = _RAND_2102[7:0];
  _RAND_2103 = {1{`RANDOM}};
  lineBuffer_2096 = _RAND_2103[7:0];
  _RAND_2104 = {1{`RANDOM}};
  lineBuffer_2097 = _RAND_2104[7:0];
  _RAND_2105 = {1{`RANDOM}};
  lineBuffer_2098 = _RAND_2105[7:0];
  _RAND_2106 = {1{`RANDOM}};
  lineBuffer_2099 = _RAND_2106[7:0];
  _RAND_2107 = {1{`RANDOM}};
  lineBuffer_2100 = _RAND_2107[7:0];
  _RAND_2108 = {1{`RANDOM}};
  lineBuffer_2101 = _RAND_2108[7:0];
  _RAND_2109 = {1{`RANDOM}};
  lineBuffer_2102 = _RAND_2109[7:0];
  _RAND_2110 = {1{`RANDOM}};
  lineBuffer_2103 = _RAND_2110[7:0];
  _RAND_2111 = {1{`RANDOM}};
  lineBuffer_2104 = _RAND_2111[7:0];
  _RAND_2112 = {1{`RANDOM}};
  lineBuffer_2105 = _RAND_2112[7:0];
  _RAND_2113 = {1{`RANDOM}};
  lineBuffer_2106 = _RAND_2113[7:0];
  _RAND_2114 = {1{`RANDOM}};
  lineBuffer_2107 = _RAND_2114[7:0];
  _RAND_2115 = {1{`RANDOM}};
  lineBuffer_2108 = _RAND_2115[7:0];
  _RAND_2116 = {1{`RANDOM}};
  lineBuffer_2109 = _RAND_2116[7:0];
  _RAND_2117 = {1{`RANDOM}};
  lineBuffer_2110 = _RAND_2117[7:0];
  _RAND_2118 = {1{`RANDOM}};
  lineBuffer_2111 = _RAND_2118[7:0];
  _RAND_2119 = {1{`RANDOM}};
  lineBuffer_2112 = _RAND_2119[7:0];
  _RAND_2120 = {1{`RANDOM}};
  lineBuffer_2113 = _RAND_2120[7:0];
  _RAND_2121 = {1{`RANDOM}};
  lineBuffer_2114 = _RAND_2121[7:0];
  _RAND_2122 = {1{`RANDOM}};
  lineBuffer_2115 = _RAND_2122[7:0];
  _RAND_2123 = {1{`RANDOM}};
  lineBuffer_2116 = _RAND_2123[7:0];
  _RAND_2124 = {1{`RANDOM}};
  lineBuffer_2117 = _RAND_2124[7:0];
  _RAND_2125 = {1{`RANDOM}};
  lineBuffer_2118 = _RAND_2125[7:0];
  _RAND_2126 = {1{`RANDOM}};
  lineBuffer_2119 = _RAND_2126[7:0];
  _RAND_2127 = {1{`RANDOM}};
  lineBuffer_2120 = _RAND_2127[7:0];
  _RAND_2128 = {1{`RANDOM}};
  lineBuffer_2121 = _RAND_2128[7:0];
  _RAND_2129 = {1{`RANDOM}};
  lineBuffer_2122 = _RAND_2129[7:0];
  _RAND_2130 = {1{`RANDOM}};
  lineBuffer_2123 = _RAND_2130[7:0];
  _RAND_2131 = {1{`RANDOM}};
  lineBuffer_2124 = _RAND_2131[7:0];
  _RAND_2132 = {1{`RANDOM}};
  lineBuffer_2125 = _RAND_2132[7:0];
  _RAND_2133 = {1{`RANDOM}};
  lineBuffer_2126 = _RAND_2133[7:0];
  _RAND_2134 = {1{`RANDOM}};
  lineBuffer_2127 = _RAND_2134[7:0];
  _RAND_2135 = {1{`RANDOM}};
  lineBuffer_2128 = _RAND_2135[7:0];
  _RAND_2136 = {1{`RANDOM}};
  lineBuffer_2129 = _RAND_2136[7:0];
  _RAND_2137 = {1{`RANDOM}};
  lineBuffer_2130 = _RAND_2137[7:0];
  _RAND_2138 = {1{`RANDOM}};
  lineBuffer_2131 = _RAND_2138[7:0];
  _RAND_2139 = {1{`RANDOM}};
  lineBuffer_2132 = _RAND_2139[7:0];
  _RAND_2140 = {1{`RANDOM}};
  lineBuffer_2133 = _RAND_2140[7:0];
  _RAND_2141 = {1{`RANDOM}};
  lineBuffer_2134 = _RAND_2141[7:0];
  _RAND_2142 = {1{`RANDOM}};
  lineBuffer_2135 = _RAND_2142[7:0];
  _RAND_2143 = {1{`RANDOM}};
  lineBuffer_2136 = _RAND_2143[7:0];
  _RAND_2144 = {1{`RANDOM}};
  lineBuffer_2137 = _RAND_2144[7:0];
  _RAND_2145 = {1{`RANDOM}};
  lineBuffer_2138 = _RAND_2145[7:0];
  _RAND_2146 = {1{`RANDOM}};
  lineBuffer_2139 = _RAND_2146[7:0];
  _RAND_2147 = {1{`RANDOM}};
  lineBuffer_2140 = _RAND_2147[7:0];
  _RAND_2148 = {1{`RANDOM}};
  lineBuffer_2141 = _RAND_2148[7:0];
  _RAND_2149 = {1{`RANDOM}};
  lineBuffer_2142 = _RAND_2149[7:0];
  _RAND_2150 = {1{`RANDOM}};
  lineBuffer_2143 = _RAND_2150[7:0];
  _RAND_2151 = {1{`RANDOM}};
  lineBuffer_2144 = _RAND_2151[7:0];
  _RAND_2152 = {1{`RANDOM}};
  lineBuffer_2145 = _RAND_2152[7:0];
  _RAND_2153 = {1{`RANDOM}};
  lineBuffer_2146 = _RAND_2153[7:0];
  _RAND_2154 = {1{`RANDOM}};
  lineBuffer_2147 = _RAND_2154[7:0];
  _RAND_2155 = {1{`RANDOM}};
  lineBuffer_2148 = _RAND_2155[7:0];
  _RAND_2156 = {1{`RANDOM}};
  lineBuffer_2149 = _RAND_2156[7:0];
  _RAND_2157 = {1{`RANDOM}};
  lineBuffer_2150 = _RAND_2157[7:0];
  _RAND_2158 = {1{`RANDOM}};
  lineBuffer_2151 = _RAND_2158[7:0];
  _RAND_2159 = {1{`RANDOM}};
  lineBuffer_2152 = _RAND_2159[7:0];
  _RAND_2160 = {1{`RANDOM}};
  lineBuffer_2153 = _RAND_2160[7:0];
  _RAND_2161 = {1{`RANDOM}};
  lineBuffer_2154 = _RAND_2161[7:0];
  _RAND_2162 = {1{`RANDOM}};
  lineBuffer_2155 = _RAND_2162[7:0];
  _RAND_2163 = {1{`RANDOM}};
  lineBuffer_2156 = _RAND_2163[7:0];
  _RAND_2164 = {1{`RANDOM}};
  lineBuffer_2157 = _RAND_2164[7:0];
  _RAND_2165 = {1{`RANDOM}};
  lineBuffer_2158 = _RAND_2165[7:0];
  _RAND_2166 = {1{`RANDOM}};
  lineBuffer_2159 = _RAND_2166[7:0];
  _RAND_2167 = {1{`RANDOM}};
  lineBuffer_2160 = _RAND_2167[7:0];
  _RAND_2168 = {1{`RANDOM}};
  lineBuffer_2161 = _RAND_2168[7:0];
  _RAND_2169 = {1{`RANDOM}};
  lineBuffer_2162 = _RAND_2169[7:0];
  _RAND_2170 = {1{`RANDOM}};
  lineBuffer_2163 = _RAND_2170[7:0];
  _RAND_2171 = {1{`RANDOM}};
  lineBuffer_2164 = _RAND_2171[7:0];
  _RAND_2172 = {1{`RANDOM}};
  lineBuffer_2165 = _RAND_2172[7:0];
  _RAND_2173 = {1{`RANDOM}};
  lineBuffer_2166 = _RAND_2173[7:0];
  _RAND_2174 = {1{`RANDOM}};
  lineBuffer_2167 = _RAND_2174[7:0];
  _RAND_2175 = {1{`RANDOM}};
  lineBuffer_2168 = _RAND_2175[7:0];
  _RAND_2176 = {1{`RANDOM}};
  lineBuffer_2169 = _RAND_2176[7:0];
  _RAND_2177 = {1{`RANDOM}};
  lineBuffer_2170 = _RAND_2177[7:0];
  _RAND_2178 = {1{`RANDOM}};
  lineBuffer_2171 = _RAND_2178[7:0];
  _RAND_2179 = {1{`RANDOM}};
  lineBuffer_2172 = _RAND_2179[7:0];
  _RAND_2180 = {1{`RANDOM}};
  lineBuffer_2173 = _RAND_2180[7:0];
  _RAND_2181 = {1{`RANDOM}};
  lineBuffer_2174 = _RAND_2181[7:0];
  _RAND_2182 = {1{`RANDOM}};
  lineBuffer_2175 = _RAND_2182[7:0];
  _RAND_2183 = {1{`RANDOM}};
  lineBuffer_2176 = _RAND_2183[7:0];
  _RAND_2184 = {1{`RANDOM}};
  lineBuffer_2177 = _RAND_2184[7:0];
  _RAND_2185 = {1{`RANDOM}};
  lineBuffer_2178 = _RAND_2185[7:0];
  _RAND_2186 = {1{`RANDOM}};
  lineBuffer_2179 = _RAND_2186[7:0];
  _RAND_2187 = {1{`RANDOM}};
  lineBuffer_2180 = _RAND_2187[7:0];
  _RAND_2188 = {1{`RANDOM}};
  lineBuffer_2181 = _RAND_2188[7:0];
  _RAND_2189 = {1{`RANDOM}};
  lineBuffer_2182 = _RAND_2189[7:0];
  _RAND_2190 = {1{`RANDOM}};
  lineBuffer_2183 = _RAND_2190[7:0];
  _RAND_2191 = {1{`RANDOM}};
  lineBuffer_2184 = _RAND_2191[7:0];
  _RAND_2192 = {1{`RANDOM}};
  lineBuffer_2185 = _RAND_2192[7:0];
  _RAND_2193 = {1{`RANDOM}};
  lineBuffer_2186 = _RAND_2193[7:0];
  _RAND_2194 = {1{`RANDOM}};
  lineBuffer_2187 = _RAND_2194[7:0];
  _RAND_2195 = {1{`RANDOM}};
  lineBuffer_2188 = _RAND_2195[7:0];
  _RAND_2196 = {1{`RANDOM}};
  lineBuffer_2189 = _RAND_2196[7:0];
  _RAND_2197 = {1{`RANDOM}};
  lineBuffer_2190 = _RAND_2197[7:0];
  _RAND_2198 = {1{`RANDOM}};
  lineBuffer_2191 = _RAND_2198[7:0];
  _RAND_2199 = {1{`RANDOM}};
  lineBuffer_2192 = _RAND_2199[7:0];
  _RAND_2200 = {1{`RANDOM}};
  lineBuffer_2193 = _RAND_2200[7:0];
  _RAND_2201 = {1{`RANDOM}};
  lineBuffer_2194 = _RAND_2201[7:0];
  _RAND_2202 = {1{`RANDOM}};
  lineBuffer_2195 = _RAND_2202[7:0];
  _RAND_2203 = {1{`RANDOM}};
  lineBuffer_2196 = _RAND_2203[7:0];
  _RAND_2204 = {1{`RANDOM}};
  lineBuffer_2197 = _RAND_2204[7:0];
  _RAND_2205 = {1{`RANDOM}};
  lineBuffer_2198 = _RAND_2205[7:0];
  _RAND_2206 = {1{`RANDOM}};
  lineBuffer_2199 = _RAND_2206[7:0];
  _RAND_2207 = {1{`RANDOM}};
  lineBuffer_2200 = _RAND_2207[7:0];
  _RAND_2208 = {1{`RANDOM}};
  lineBuffer_2201 = _RAND_2208[7:0];
  _RAND_2209 = {1{`RANDOM}};
  lineBuffer_2202 = _RAND_2209[7:0];
  _RAND_2210 = {1{`RANDOM}};
  lineBuffer_2203 = _RAND_2210[7:0];
  _RAND_2211 = {1{`RANDOM}};
  lineBuffer_2204 = _RAND_2211[7:0];
  _RAND_2212 = {1{`RANDOM}};
  lineBuffer_2205 = _RAND_2212[7:0];
  _RAND_2213 = {1{`RANDOM}};
  lineBuffer_2206 = _RAND_2213[7:0];
  _RAND_2214 = {1{`RANDOM}};
  lineBuffer_2207 = _RAND_2214[7:0];
  _RAND_2215 = {1{`RANDOM}};
  lineBuffer_2208 = _RAND_2215[7:0];
  _RAND_2216 = {1{`RANDOM}};
  lineBuffer_2209 = _RAND_2216[7:0];
  _RAND_2217 = {1{`RANDOM}};
  lineBuffer_2210 = _RAND_2217[7:0];
  _RAND_2218 = {1{`RANDOM}};
  lineBuffer_2211 = _RAND_2218[7:0];
  _RAND_2219 = {1{`RANDOM}};
  lineBuffer_2212 = _RAND_2219[7:0];
  _RAND_2220 = {1{`RANDOM}};
  lineBuffer_2213 = _RAND_2220[7:0];
  _RAND_2221 = {1{`RANDOM}};
  lineBuffer_2214 = _RAND_2221[7:0];
  _RAND_2222 = {1{`RANDOM}};
  lineBuffer_2215 = _RAND_2222[7:0];
  _RAND_2223 = {1{`RANDOM}};
  lineBuffer_2216 = _RAND_2223[7:0];
  _RAND_2224 = {1{`RANDOM}};
  lineBuffer_2217 = _RAND_2224[7:0];
  _RAND_2225 = {1{`RANDOM}};
  lineBuffer_2218 = _RAND_2225[7:0];
  _RAND_2226 = {1{`RANDOM}};
  lineBuffer_2219 = _RAND_2226[7:0];
  _RAND_2227 = {1{`RANDOM}};
  lineBuffer_2220 = _RAND_2227[7:0];
  _RAND_2228 = {1{`RANDOM}};
  lineBuffer_2221 = _RAND_2228[7:0];
  _RAND_2229 = {1{`RANDOM}};
  lineBuffer_2222 = _RAND_2229[7:0];
  _RAND_2230 = {1{`RANDOM}};
  lineBuffer_2223 = _RAND_2230[7:0];
  _RAND_2231 = {1{`RANDOM}};
  lineBuffer_2224 = _RAND_2231[7:0];
  _RAND_2232 = {1{`RANDOM}};
  lineBuffer_2225 = _RAND_2232[7:0];
  _RAND_2233 = {1{`RANDOM}};
  lineBuffer_2226 = _RAND_2233[7:0];
  _RAND_2234 = {1{`RANDOM}};
  lineBuffer_2227 = _RAND_2234[7:0];
  _RAND_2235 = {1{`RANDOM}};
  lineBuffer_2228 = _RAND_2235[7:0];
  _RAND_2236 = {1{`RANDOM}};
  lineBuffer_2229 = _RAND_2236[7:0];
  _RAND_2237 = {1{`RANDOM}};
  lineBuffer_2230 = _RAND_2237[7:0];
  _RAND_2238 = {1{`RANDOM}};
  lineBuffer_2231 = _RAND_2238[7:0];
  _RAND_2239 = {1{`RANDOM}};
  lineBuffer_2232 = _RAND_2239[7:0];
  _RAND_2240 = {1{`RANDOM}};
  lineBuffer_2233 = _RAND_2240[7:0];
  _RAND_2241 = {1{`RANDOM}};
  lineBuffer_2234 = _RAND_2241[7:0];
  _RAND_2242 = {1{`RANDOM}};
  lineBuffer_2235 = _RAND_2242[7:0];
  _RAND_2243 = {1{`RANDOM}};
  lineBuffer_2236 = _RAND_2243[7:0];
  _RAND_2244 = {1{`RANDOM}};
  lineBuffer_2237 = _RAND_2244[7:0];
  _RAND_2245 = {1{`RANDOM}};
  lineBuffer_2238 = _RAND_2245[7:0];
  _RAND_2246 = {1{`RANDOM}};
  lineBuffer_2239 = _RAND_2246[7:0];
  _RAND_2247 = {1{`RANDOM}};
  lineBuffer_2240 = _RAND_2247[7:0];
  _RAND_2248 = {1{`RANDOM}};
  lineBuffer_2241 = _RAND_2248[7:0];
  _RAND_2249 = {1{`RANDOM}};
  lineBuffer_2242 = _RAND_2249[7:0];
  _RAND_2250 = {1{`RANDOM}};
  lineBuffer_2243 = _RAND_2250[7:0];
  _RAND_2251 = {1{`RANDOM}};
  lineBuffer_2244 = _RAND_2251[7:0];
  _RAND_2252 = {1{`RANDOM}};
  lineBuffer_2245 = _RAND_2252[7:0];
  _RAND_2253 = {1{`RANDOM}};
  lineBuffer_2246 = _RAND_2253[7:0];
  _RAND_2254 = {1{`RANDOM}};
  lineBuffer_2247 = _RAND_2254[7:0];
  _RAND_2255 = {1{`RANDOM}};
  lineBuffer_2248 = _RAND_2255[7:0];
  _RAND_2256 = {1{`RANDOM}};
  lineBuffer_2249 = _RAND_2256[7:0];
  _RAND_2257 = {1{`RANDOM}};
  lineBuffer_2250 = _RAND_2257[7:0];
  _RAND_2258 = {1{`RANDOM}};
  lineBuffer_2251 = _RAND_2258[7:0];
  _RAND_2259 = {1{`RANDOM}};
  lineBuffer_2252 = _RAND_2259[7:0];
  _RAND_2260 = {1{`RANDOM}};
  lineBuffer_2253 = _RAND_2260[7:0];
  _RAND_2261 = {1{`RANDOM}};
  lineBuffer_2254 = _RAND_2261[7:0];
  _RAND_2262 = {1{`RANDOM}};
  lineBuffer_2255 = _RAND_2262[7:0];
  _RAND_2263 = {1{`RANDOM}};
  lineBuffer_2256 = _RAND_2263[7:0];
  _RAND_2264 = {1{`RANDOM}};
  lineBuffer_2257 = _RAND_2264[7:0];
  _RAND_2265 = {1{`RANDOM}};
  lineBuffer_2258 = _RAND_2265[7:0];
  _RAND_2266 = {1{`RANDOM}};
  lineBuffer_2259 = _RAND_2266[7:0];
  _RAND_2267 = {1{`RANDOM}};
  lineBuffer_2260 = _RAND_2267[7:0];
  _RAND_2268 = {1{`RANDOM}};
  lineBuffer_2261 = _RAND_2268[7:0];
  _RAND_2269 = {1{`RANDOM}};
  lineBuffer_2262 = _RAND_2269[7:0];
  _RAND_2270 = {1{`RANDOM}};
  lineBuffer_2263 = _RAND_2270[7:0];
  _RAND_2271 = {1{`RANDOM}};
  lineBuffer_2264 = _RAND_2271[7:0];
  _RAND_2272 = {1{`RANDOM}};
  lineBuffer_2265 = _RAND_2272[7:0];
  _RAND_2273 = {1{`RANDOM}};
  lineBuffer_2266 = _RAND_2273[7:0];
  _RAND_2274 = {1{`RANDOM}};
  lineBuffer_2267 = _RAND_2274[7:0];
  _RAND_2275 = {1{`RANDOM}};
  lineBuffer_2268 = _RAND_2275[7:0];
  _RAND_2276 = {1{`RANDOM}};
  lineBuffer_2269 = _RAND_2276[7:0];
  _RAND_2277 = {1{`RANDOM}};
  lineBuffer_2270 = _RAND_2277[7:0];
  _RAND_2278 = {1{`RANDOM}};
  lineBuffer_2271 = _RAND_2278[7:0];
  _RAND_2279 = {1{`RANDOM}};
  lineBuffer_2272 = _RAND_2279[7:0];
  _RAND_2280 = {1{`RANDOM}};
  lineBuffer_2273 = _RAND_2280[7:0];
  _RAND_2281 = {1{`RANDOM}};
  lineBuffer_2274 = _RAND_2281[7:0];
  _RAND_2282 = {1{`RANDOM}};
  lineBuffer_2275 = _RAND_2282[7:0];
  _RAND_2283 = {1{`RANDOM}};
  lineBuffer_2276 = _RAND_2283[7:0];
  _RAND_2284 = {1{`RANDOM}};
  lineBuffer_2277 = _RAND_2284[7:0];
  _RAND_2285 = {1{`RANDOM}};
  lineBuffer_2278 = _RAND_2285[7:0];
  _RAND_2286 = {1{`RANDOM}};
  lineBuffer_2279 = _RAND_2286[7:0];
  _RAND_2287 = {1{`RANDOM}};
  lineBuffer_2280 = _RAND_2287[7:0];
  _RAND_2288 = {1{`RANDOM}};
  lineBuffer_2281 = _RAND_2288[7:0];
  _RAND_2289 = {1{`RANDOM}};
  lineBuffer_2282 = _RAND_2289[7:0];
  _RAND_2290 = {1{`RANDOM}};
  lineBuffer_2283 = _RAND_2290[7:0];
  _RAND_2291 = {1{`RANDOM}};
  lineBuffer_2284 = _RAND_2291[7:0];
  _RAND_2292 = {1{`RANDOM}};
  lineBuffer_2285 = _RAND_2292[7:0];
  _RAND_2293 = {1{`RANDOM}};
  lineBuffer_2286 = _RAND_2293[7:0];
  _RAND_2294 = {1{`RANDOM}};
  lineBuffer_2287 = _RAND_2294[7:0];
  _RAND_2295 = {1{`RANDOM}};
  lineBuffer_2288 = _RAND_2295[7:0];
  _RAND_2296 = {1{`RANDOM}};
  lineBuffer_2289 = _RAND_2296[7:0];
  _RAND_2297 = {1{`RANDOM}};
  lineBuffer_2290 = _RAND_2297[7:0];
  _RAND_2298 = {1{`RANDOM}};
  lineBuffer_2291 = _RAND_2298[7:0];
  _RAND_2299 = {1{`RANDOM}};
  lineBuffer_2292 = _RAND_2299[7:0];
  _RAND_2300 = {1{`RANDOM}};
  lineBuffer_2293 = _RAND_2300[7:0];
  _RAND_2301 = {1{`RANDOM}};
  lineBuffer_2294 = _RAND_2301[7:0];
  _RAND_2302 = {1{`RANDOM}};
  lineBuffer_2295 = _RAND_2302[7:0];
  _RAND_2303 = {1{`RANDOM}};
  lineBuffer_2296 = _RAND_2303[7:0];
  _RAND_2304 = {1{`RANDOM}};
  lineBuffer_2297 = _RAND_2304[7:0];
  _RAND_2305 = {1{`RANDOM}};
  lineBuffer_2298 = _RAND_2305[7:0];
  _RAND_2306 = {1{`RANDOM}};
  lineBuffer_2299 = _RAND_2306[7:0];
  _RAND_2307 = {1{`RANDOM}};
  lineBuffer_2300 = _RAND_2307[7:0];
  _RAND_2308 = {1{`RANDOM}};
  lineBuffer_2301 = _RAND_2308[7:0];
  _RAND_2309 = {1{`RANDOM}};
  lineBuffer_2302 = _RAND_2309[7:0];
  _RAND_2310 = {1{`RANDOM}};
  lineBuffer_2303 = _RAND_2310[7:0];
  _RAND_2311 = {1{`RANDOM}};
  lineBuffer_2304 = _RAND_2311[7:0];
  _RAND_2312 = {1{`RANDOM}};
  lineBuffer_2305 = _RAND_2312[7:0];
  _RAND_2313 = {1{`RANDOM}};
  lineBuffer_2306 = _RAND_2313[7:0];
  _RAND_2314 = {1{`RANDOM}};
  lineBuffer_2307 = _RAND_2314[7:0];
  _RAND_2315 = {1{`RANDOM}};
  lineBuffer_2308 = _RAND_2315[7:0];
  _RAND_2316 = {1{`RANDOM}};
  lineBuffer_2309 = _RAND_2316[7:0];
  _RAND_2317 = {1{`RANDOM}};
  lineBuffer_2310 = _RAND_2317[7:0];
  _RAND_2318 = {1{`RANDOM}};
  lineBuffer_2311 = _RAND_2318[7:0];
  _RAND_2319 = {1{`RANDOM}};
  lineBuffer_2312 = _RAND_2319[7:0];
  _RAND_2320 = {1{`RANDOM}};
  lineBuffer_2313 = _RAND_2320[7:0];
  _RAND_2321 = {1{`RANDOM}};
  lineBuffer_2314 = _RAND_2321[7:0];
  _RAND_2322 = {1{`RANDOM}};
  lineBuffer_2315 = _RAND_2322[7:0];
  _RAND_2323 = {1{`RANDOM}};
  lineBuffer_2316 = _RAND_2323[7:0];
  _RAND_2324 = {1{`RANDOM}};
  lineBuffer_2317 = _RAND_2324[7:0];
  _RAND_2325 = {1{`RANDOM}};
  lineBuffer_2318 = _RAND_2325[7:0];
  _RAND_2326 = {1{`RANDOM}};
  lineBuffer_2319 = _RAND_2326[7:0];
  _RAND_2327 = {1{`RANDOM}};
  lineBuffer_2320 = _RAND_2327[7:0];
  _RAND_2328 = {1{`RANDOM}};
  lineBuffer_2321 = _RAND_2328[7:0];
  _RAND_2329 = {1{`RANDOM}};
  lineBuffer_2322 = _RAND_2329[7:0];
  _RAND_2330 = {1{`RANDOM}};
  lineBuffer_2323 = _RAND_2330[7:0];
  _RAND_2331 = {1{`RANDOM}};
  lineBuffer_2324 = _RAND_2331[7:0];
  _RAND_2332 = {1{`RANDOM}};
  lineBuffer_2325 = _RAND_2332[7:0];
  _RAND_2333 = {1{`RANDOM}};
  lineBuffer_2326 = _RAND_2333[7:0];
  _RAND_2334 = {1{`RANDOM}};
  lineBuffer_2327 = _RAND_2334[7:0];
  _RAND_2335 = {1{`RANDOM}};
  lineBuffer_2328 = _RAND_2335[7:0];
  _RAND_2336 = {1{`RANDOM}};
  lineBuffer_2329 = _RAND_2336[7:0];
  _RAND_2337 = {1{`RANDOM}};
  lineBuffer_2330 = _RAND_2337[7:0];
  _RAND_2338 = {1{`RANDOM}};
  lineBuffer_2331 = _RAND_2338[7:0];
  _RAND_2339 = {1{`RANDOM}};
  lineBuffer_2332 = _RAND_2339[7:0];
  _RAND_2340 = {1{`RANDOM}};
  lineBuffer_2333 = _RAND_2340[7:0];
  _RAND_2341 = {1{`RANDOM}};
  lineBuffer_2334 = _RAND_2341[7:0];
  _RAND_2342 = {1{`RANDOM}};
  lineBuffer_2335 = _RAND_2342[7:0];
  _RAND_2343 = {1{`RANDOM}};
  lineBuffer_2336 = _RAND_2343[7:0];
  _RAND_2344 = {1{`RANDOM}};
  lineBuffer_2337 = _RAND_2344[7:0];
  _RAND_2345 = {1{`RANDOM}};
  lineBuffer_2338 = _RAND_2345[7:0];
  _RAND_2346 = {1{`RANDOM}};
  lineBuffer_2339 = _RAND_2346[7:0];
  _RAND_2347 = {1{`RANDOM}};
  lineBuffer_2340 = _RAND_2347[7:0];
  _RAND_2348 = {1{`RANDOM}};
  lineBuffer_2341 = _RAND_2348[7:0];
  _RAND_2349 = {1{`RANDOM}};
  lineBuffer_2342 = _RAND_2349[7:0];
  _RAND_2350 = {1{`RANDOM}};
  lineBuffer_2343 = _RAND_2350[7:0];
  _RAND_2351 = {1{`RANDOM}};
  lineBuffer_2344 = _RAND_2351[7:0];
  _RAND_2352 = {1{`RANDOM}};
  lineBuffer_2345 = _RAND_2352[7:0];
  _RAND_2353 = {1{`RANDOM}};
  lineBuffer_2346 = _RAND_2353[7:0];
  _RAND_2354 = {1{`RANDOM}};
  lineBuffer_2347 = _RAND_2354[7:0];
  _RAND_2355 = {1{`RANDOM}};
  lineBuffer_2348 = _RAND_2355[7:0];
  _RAND_2356 = {1{`RANDOM}};
  lineBuffer_2349 = _RAND_2356[7:0];
  _RAND_2357 = {1{`RANDOM}};
  lineBuffer_2350 = _RAND_2357[7:0];
  _RAND_2358 = {1{`RANDOM}};
  lineBuffer_2351 = _RAND_2358[7:0];
  _RAND_2359 = {1{`RANDOM}};
  lineBuffer_2352 = _RAND_2359[7:0];
  _RAND_2360 = {1{`RANDOM}};
  lineBuffer_2353 = _RAND_2360[7:0];
  _RAND_2361 = {1{`RANDOM}};
  lineBuffer_2354 = _RAND_2361[7:0];
  _RAND_2362 = {1{`RANDOM}};
  lineBuffer_2355 = _RAND_2362[7:0];
  _RAND_2363 = {1{`RANDOM}};
  lineBuffer_2356 = _RAND_2363[7:0];
  _RAND_2364 = {1{`RANDOM}};
  lineBuffer_2357 = _RAND_2364[7:0];
  _RAND_2365 = {1{`RANDOM}};
  lineBuffer_2358 = _RAND_2365[7:0];
  _RAND_2366 = {1{`RANDOM}};
  lineBuffer_2359 = _RAND_2366[7:0];
  _RAND_2367 = {1{`RANDOM}};
  lineBuffer_2360 = _RAND_2367[7:0];
  _RAND_2368 = {1{`RANDOM}};
  lineBuffer_2361 = _RAND_2368[7:0];
  _RAND_2369 = {1{`RANDOM}};
  lineBuffer_2362 = _RAND_2369[7:0];
  _RAND_2370 = {1{`RANDOM}};
  lineBuffer_2363 = _RAND_2370[7:0];
  _RAND_2371 = {1{`RANDOM}};
  lineBuffer_2364 = _RAND_2371[7:0];
  _RAND_2372 = {1{`RANDOM}};
  lineBuffer_2365 = _RAND_2372[7:0];
  _RAND_2373 = {1{`RANDOM}};
  lineBuffer_2366 = _RAND_2373[7:0];
  _RAND_2374 = {1{`RANDOM}};
  lineBuffer_2367 = _RAND_2374[7:0];
  _RAND_2375 = {1{`RANDOM}};
  lineBuffer_2368 = _RAND_2375[7:0];
  _RAND_2376 = {1{`RANDOM}};
  lineBuffer_2369 = _RAND_2376[7:0];
  _RAND_2377 = {1{`RANDOM}};
  lineBuffer_2370 = _RAND_2377[7:0];
  _RAND_2378 = {1{`RANDOM}};
  lineBuffer_2371 = _RAND_2378[7:0];
  _RAND_2379 = {1{`RANDOM}};
  lineBuffer_2372 = _RAND_2379[7:0];
  _RAND_2380 = {1{`RANDOM}};
  lineBuffer_2373 = _RAND_2380[7:0];
  _RAND_2381 = {1{`RANDOM}};
  lineBuffer_2374 = _RAND_2381[7:0];
  _RAND_2382 = {1{`RANDOM}};
  lineBuffer_2375 = _RAND_2382[7:0];
  _RAND_2383 = {1{`RANDOM}};
  lineBuffer_2376 = _RAND_2383[7:0];
  _RAND_2384 = {1{`RANDOM}};
  lineBuffer_2377 = _RAND_2384[7:0];
  _RAND_2385 = {1{`RANDOM}};
  lineBuffer_2378 = _RAND_2385[7:0];
  _RAND_2386 = {1{`RANDOM}};
  lineBuffer_2379 = _RAND_2386[7:0];
  _RAND_2387 = {1{`RANDOM}};
  lineBuffer_2380 = _RAND_2387[7:0];
  _RAND_2388 = {1{`RANDOM}};
  lineBuffer_2381 = _RAND_2388[7:0];
  _RAND_2389 = {1{`RANDOM}};
  lineBuffer_2382 = _RAND_2389[7:0];
  _RAND_2390 = {1{`RANDOM}};
  lineBuffer_2383 = _RAND_2390[7:0];
  _RAND_2391 = {1{`RANDOM}};
  lineBuffer_2384 = _RAND_2391[7:0];
  _RAND_2392 = {1{`RANDOM}};
  lineBuffer_2385 = _RAND_2392[7:0];
  _RAND_2393 = {1{`RANDOM}};
  lineBuffer_2386 = _RAND_2393[7:0];
  _RAND_2394 = {1{`RANDOM}};
  lineBuffer_2387 = _RAND_2394[7:0];
  _RAND_2395 = {1{`RANDOM}};
  lineBuffer_2388 = _RAND_2395[7:0];
  _RAND_2396 = {1{`RANDOM}};
  lineBuffer_2389 = _RAND_2396[7:0];
  _RAND_2397 = {1{`RANDOM}};
  lineBuffer_2390 = _RAND_2397[7:0];
  _RAND_2398 = {1{`RANDOM}};
  lineBuffer_2391 = _RAND_2398[7:0];
  _RAND_2399 = {1{`RANDOM}};
  lineBuffer_2392 = _RAND_2399[7:0];
  _RAND_2400 = {1{`RANDOM}};
  lineBuffer_2393 = _RAND_2400[7:0];
  _RAND_2401 = {1{`RANDOM}};
  lineBuffer_2394 = _RAND_2401[7:0];
  _RAND_2402 = {1{`RANDOM}};
  lineBuffer_2395 = _RAND_2402[7:0];
  _RAND_2403 = {1{`RANDOM}};
  lineBuffer_2396 = _RAND_2403[7:0];
  _RAND_2404 = {1{`RANDOM}};
  lineBuffer_2397 = _RAND_2404[7:0];
  _RAND_2405 = {1{`RANDOM}};
  lineBuffer_2398 = _RAND_2405[7:0];
  _RAND_2406 = {1{`RANDOM}};
  lineBuffer_2399 = _RAND_2406[7:0];
  _RAND_2407 = {1{`RANDOM}};
  lineBuffer_2400 = _RAND_2407[7:0];
  _RAND_2408 = {1{`RANDOM}};
  lineBuffer_2401 = _RAND_2408[7:0];
  _RAND_2409 = {1{`RANDOM}};
  lineBuffer_2402 = _RAND_2409[7:0];
  _RAND_2410 = {1{`RANDOM}};
  lineBuffer_2403 = _RAND_2410[7:0];
  _RAND_2411 = {1{`RANDOM}};
  lineBuffer_2404 = _RAND_2411[7:0];
  _RAND_2412 = {1{`RANDOM}};
  lineBuffer_2405 = _RAND_2412[7:0];
  _RAND_2413 = {1{`RANDOM}};
  lineBuffer_2406 = _RAND_2413[7:0];
  _RAND_2414 = {1{`RANDOM}};
  lineBuffer_2407 = _RAND_2414[7:0];
  _RAND_2415 = {1{`RANDOM}};
  lineBuffer_2408 = _RAND_2415[7:0];
  _RAND_2416 = {1{`RANDOM}};
  lineBuffer_2409 = _RAND_2416[7:0];
  _RAND_2417 = {1{`RANDOM}};
  lineBuffer_2410 = _RAND_2417[7:0];
  _RAND_2418 = {1{`RANDOM}};
  lineBuffer_2411 = _RAND_2418[7:0];
  _RAND_2419 = {1{`RANDOM}};
  lineBuffer_2412 = _RAND_2419[7:0];
  _RAND_2420 = {1{`RANDOM}};
  lineBuffer_2413 = _RAND_2420[7:0];
  _RAND_2421 = {1{`RANDOM}};
  lineBuffer_2414 = _RAND_2421[7:0];
  _RAND_2422 = {1{`RANDOM}};
  lineBuffer_2415 = _RAND_2422[7:0];
  _RAND_2423 = {1{`RANDOM}};
  lineBuffer_2416 = _RAND_2423[7:0];
  _RAND_2424 = {1{`RANDOM}};
  lineBuffer_2417 = _RAND_2424[7:0];
  _RAND_2425 = {1{`RANDOM}};
  lineBuffer_2418 = _RAND_2425[7:0];
  _RAND_2426 = {1{`RANDOM}};
  lineBuffer_2419 = _RAND_2426[7:0];
  _RAND_2427 = {1{`RANDOM}};
  lineBuffer_2420 = _RAND_2427[7:0];
  _RAND_2428 = {1{`RANDOM}};
  lineBuffer_2421 = _RAND_2428[7:0];
  _RAND_2429 = {1{`RANDOM}};
  lineBuffer_2422 = _RAND_2429[7:0];
  _RAND_2430 = {1{`RANDOM}};
  lineBuffer_2423 = _RAND_2430[7:0];
  _RAND_2431 = {1{`RANDOM}};
  lineBuffer_2424 = _RAND_2431[7:0];
  _RAND_2432 = {1{`RANDOM}};
  lineBuffer_2425 = _RAND_2432[7:0];
  _RAND_2433 = {1{`RANDOM}};
  lineBuffer_2426 = _RAND_2433[7:0];
  _RAND_2434 = {1{`RANDOM}};
  lineBuffer_2427 = _RAND_2434[7:0];
  _RAND_2435 = {1{`RANDOM}};
  lineBuffer_2428 = _RAND_2435[7:0];
  _RAND_2436 = {1{`RANDOM}};
  lineBuffer_2429 = _RAND_2436[7:0];
  _RAND_2437 = {1{`RANDOM}};
  lineBuffer_2430 = _RAND_2437[7:0];
  _RAND_2438 = {1{`RANDOM}};
  lineBuffer_2431 = _RAND_2438[7:0];
  _RAND_2439 = {1{`RANDOM}};
  lineBuffer_2432 = _RAND_2439[7:0];
  _RAND_2440 = {1{`RANDOM}};
  lineBuffer_2433 = _RAND_2440[7:0];
  _RAND_2441 = {1{`RANDOM}};
  lineBuffer_2434 = _RAND_2441[7:0];
  _RAND_2442 = {1{`RANDOM}};
  lineBuffer_2435 = _RAND_2442[7:0];
  _RAND_2443 = {1{`RANDOM}};
  lineBuffer_2436 = _RAND_2443[7:0];
  _RAND_2444 = {1{`RANDOM}};
  lineBuffer_2437 = _RAND_2444[7:0];
  _RAND_2445 = {1{`RANDOM}};
  lineBuffer_2438 = _RAND_2445[7:0];
  _RAND_2446 = {1{`RANDOM}};
  lineBuffer_2439 = _RAND_2446[7:0];
  _RAND_2447 = {1{`RANDOM}};
  lineBuffer_2440 = _RAND_2447[7:0];
  _RAND_2448 = {1{`RANDOM}};
  lineBuffer_2441 = _RAND_2448[7:0];
  _RAND_2449 = {1{`RANDOM}};
  lineBuffer_2442 = _RAND_2449[7:0];
  _RAND_2450 = {1{`RANDOM}};
  lineBuffer_2443 = _RAND_2450[7:0];
  _RAND_2451 = {1{`RANDOM}};
  lineBuffer_2444 = _RAND_2451[7:0];
  _RAND_2452 = {1{`RANDOM}};
  lineBuffer_2445 = _RAND_2452[7:0];
  _RAND_2453 = {1{`RANDOM}};
  lineBuffer_2446 = _RAND_2453[7:0];
  _RAND_2454 = {1{`RANDOM}};
  lineBuffer_2447 = _RAND_2454[7:0];
  _RAND_2455 = {1{`RANDOM}};
  lineBuffer_2448 = _RAND_2455[7:0];
  _RAND_2456 = {1{`RANDOM}};
  lineBuffer_2449 = _RAND_2456[7:0];
  _RAND_2457 = {1{`RANDOM}};
  lineBuffer_2450 = _RAND_2457[7:0];
  _RAND_2458 = {1{`RANDOM}};
  lineBuffer_2451 = _RAND_2458[7:0];
  _RAND_2459 = {1{`RANDOM}};
  lineBuffer_2452 = _RAND_2459[7:0];
  _RAND_2460 = {1{`RANDOM}};
  lineBuffer_2453 = _RAND_2460[7:0];
  _RAND_2461 = {1{`RANDOM}};
  lineBuffer_2454 = _RAND_2461[7:0];
  _RAND_2462 = {1{`RANDOM}};
  lineBuffer_2455 = _RAND_2462[7:0];
  _RAND_2463 = {1{`RANDOM}};
  lineBuffer_2456 = _RAND_2463[7:0];
  _RAND_2464 = {1{`RANDOM}};
  lineBuffer_2457 = _RAND_2464[7:0];
  _RAND_2465 = {1{`RANDOM}};
  lineBuffer_2458 = _RAND_2465[7:0];
  _RAND_2466 = {1{`RANDOM}};
  lineBuffer_2459 = _RAND_2466[7:0];
  _RAND_2467 = {1{`RANDOM}};
  lineBuffer_2460 = _RAND_2467[7:0];
  _RAND_2468 = {1{`RANDOM}};
  lineBuffer_2461 = _RAND_2468[7:0];
  _RAND_2469 = {1{`RANDOM}};
  lineBuffer_2462 = _RAND_2469[7:0];
  _RAND_2470 = {1{`RANDOM}};
  lineBuffer_2463 = _RAND_2470[7:0];
  _RAND_2471 = {1{`RANDOM}};
  lineBuffer_2464 = _RAND_2471[7:0];
  _RAND_2472 = {1{`RANDOM}};
  lineBuffer_2465 = _RAND_2472[7:0];
  _RAND_2473 = {1{`RANDOM}};
  lineBuffer_2466 = _RAND_2473[7:0];
  _RAND_2474 = {1{`RANDOM}};
  lineBuffer_2467 = _RAND_2474[7:0];
  _RAND_2475 = {1{`RANDOM}};
  lineBuffer_2468 = _RAND_2475[7:0];
  _RAND_2476 = {1{`RANDOM}};
  lineBuffer_2469 = _RAND_2476[7:0];
  _RAND_2477 = {1{`RANDOM}};
  lineBuffer_2470 = _RAND_2477[7:0];
  _RAND_2478 = {1{`RANDOM}};
  lineBuffer_2471 = _RAND_2478[7:0];
  _RAND_2479 = {1{`RANDOM}};
  lineBuffer_2472 = _RAND_2479[7:0];
  _RAND_2480 = {1{`RANDOM}};
  lineBuffer_2473 = _RAND_2480[7:0];
  _RAND_2481 = {1{`RANDOM}};
  lineBuffer_2474 = _RAND_2481[7:0];
  _RAND_2482 = {1{`RANDOM}};
  lineBuffer_2475 = _RAND_2482[7:0];
  _RAND_2483 = {1{`RANDOM}};
  lineBuffer_2476 = _RAND_2483[7:0];
  _RAND_2484 = {1{`RANDOM}};
  lineBuffer_2477 = _RAND_2484[7:0];
  _RAND_2485 = {1{`RANDOM}};
  lineBuffer_2478 = _RAND_2485[7:0];
  _RAND_2486 = {1{`RANDOM}};
  lineBuffer_2479 = _RAND_2486[7:0];
  _RAND_2487 = {1{`RANDOM}};
  lineBuffer_2480 = _RAND_2487[7:0];
  _RAND_2488 = {1{`RANDOM}};
  lineBuffer_2481 = _RAND_2488[7:0];
  _RAND_2489 = {1{`RANDOM}};
  lineBuffer_2482 = _RAND_2489[7:0];
  _RAND_2490 = {1{`RANDOM}};
  lineBuffer_2483 = _RAND_2490[7:0];
  _RAND_2491 = {1{`RANDOM}};
  lineBuffer_2484 = _RAND_2491[7:0];
  _RAND_2492 = {1{`RANDOM}};
  lineBuffer_2485 = _RAND_2492[7:0];
  _RAND_2493 = {1{`RANDOM}};
  lineBuffer_2486 = _RAND_2493[7:0];
  _RAND_2494 = {1{`RANDOM}};
  lineBuffer_2487 = _RAND_2494[7:0];
  _RAND_2495 = {1{`RANDOM}};
  lineBuffer_2488 = _RAND_2495[7:0];
  _RAND_2496 = {1{`RANDOM}};
  lineBuffer_2489 = _RAND_2496[7:0];
  _RAND_2497 = {1{`RANDOM}};
  lineBuffer_2490 = _RAND_2497[7:0];
  _RAND_2498 = {1{`RANDOM}};
  lineBuffer_2491 = _RAND_2498[7:0];
  _RAND_2499 = {1{`RANDOM}};
  lineBuffer_2492 = _RAND_2499[7:0];
  _RAND_2500 = {1{`RANDOM}};
  lineBuffer_2493 = _RAND_2500[7:0];
  _RAND_2501 = {1{`RANDOM}};
  lineBuffer_2494 = _RAND_2501[7:0];
  _RAND_2502 = {1{`RANDOM}};
  lineBuffer_2495 = _RAND_2502[7:0];
  _RAND_2503 = {1{`RANDOM}};
  lineBuffer_2496 = _RAND_2503[7:0];
  _RAND_2504 = {1{`RANDOM}};
  lineBuffer_2497 = _RAND_2504[7:0];
  _RAND_2505 = {1{`RANDOM}};
  lineBuffer_2498 = _RAND_2505[7:0];
  _RAND_2506 = {1{`RANDOM}};
  lineBuffer_2499 = _RAND_2506[7:0];
  _RAND_2507 = {1{`RANDOM}};
  lineBuffer_2500 = _RAND_2507[7:0];
  _RAND_2508 = {1{`RANDOM}};
  lineBuffer_2501 = _RAND_2508[7:0];
  _RAND_2509 = {1{`RANDOM}};
  lineBuffer_2502 = _RAND_2509[7:0];
  _RAND_2510 = {1{`RANDOM}};
  lineBuffer_2503 = _RAND_2510[7:0];
  _RAND_2511 = {1{`RANDOM}};
  lineBuffer_2504 = _RAND_2511[7:0];
  _RAND_2512 = {1{`RANDOM}};
  lineBuffer_2505 = _RAND_2512[7:0];
  _RAND_2513 = {1{`RANDOM}};
  lineBuffer_2506 = _RAND_2513[7:0];
  _RAND_2514 = {1{`RANDOM}};
  lineBuffer_2507 = _RAND_2514[7:0];
  _RAND_2515 = {1{`RANDOM}};
  lineBuffer_2508 = _RAND_2515[7:0];
  _RAND_2516 = {1{`RANDOM}};
  lineBuffer_2509 = _RAND_2516[7:0];
  _RAND_2517 = {1{`RANDOM}};
  lineBuffer_2510 = _RAND_2517[7:0];
  _RAND_2518 = {1{`RANDOM}};
  lineBuffer_2511 = _RAND_2518[7:0];
  _RAND_2519 = {1{`RANDOM}};
  lineBuffer_2512 = _RAND_2519[7:0];
  _RAND_2520 = {1{`RANDOM}};
  lineBuffer_2513 = _RAND_2520[7:0];
  _RAND_2521 = {1{`RANDOM}};
  lineBuffer_2514 = _RAND_2521[7:0];
  _RAND_2522 = {1{`RANDOM}};
  lineBuffer_2515 = _RAND_2522[7:0];
  _RAND_2523 = {1{`RANDOM}};
  lineBuffer_2516 = _RAND_2523[7:0];
  _RAND_2524 = {1{`RANDOM}};
  lineBuffer_2517 = _RAND_2524[7:0];
  _RAND_2525 = {1{`RANDOM}};
  lineBuffer_2518 = _RAND_2525[7:0];
  _RAND_2526 = {1{`RANDOM}};
  lineBuffer_2519 = _RAND_2526[7:0];
  _RAND_2527 = {1{`RANDOM}};
  lineBuffer_2520 = _RAND_2527[7:0];
  _RAND_2528 = {1{`RANDOM}};
  lineBuffer_2521 = _RAND_2528[7:0];
  _RAND_2529 = {1{`RANDOM}};
  lineBuffer_2522 = _RAND_2529[7:0];
  _RAND_2530 = {1{`RANDOM}};
  lineBuffer_2523 = _RAND_2530[7:0];
  _RAND_2531 = {1{`RANDOM}};
  lineBuffer_2524 = _RAND_2531[7:0];
  _RAND_2532 = {1{`RANDOM}};
  lineBuffer_2525 = _RAND_2532[7:0];
  _RAND_2533 = {1{`RANDOM}};
  lineBuffer_2526 = _RAND_2533[7:0];
  _RAND_2534 = {1{`RANDOM}};
  lineBuffer_2527 = _RAND_2534[7:0];
  _RAND_2535 = {1{`RANDOM}};
  lineBuffer_2528 = _RAND_2535[7:0];
  _RAND_2536 = {1{`RANDOM}};
  lineBuffer_2529 = _RAND_2536[7:0];
  _RAND_2537 = {1{`RANDOM}};
  lineBuffer_2530 = _RAND_2537[7:0];
  _RAND_2538 = {1{`RANDOM}};
  lineBuffer_2531 = _RAND_2538[7:0];
  _RAND_2539 = {1{`RANDOM}};
  lineBuffer_2532 = _RAND_2539[7:0];
  _RAND_2540 = {1{`RANDOM}};
  lineBuffer_2533 = _RAND_2540[7:0];
  _RAND_2541 = {1{`RANDOM}};
  lineBuffer_2534 = _RAND_2541[7:0];
  _RAND_2542 = {1{`RANDOM}};
  lineBuffer_2535 = _RAND_2542[7:0];
  _RAND_2543 = {1{`RANDOM}};
  lineBuffer_2536 = _RAND_2543[7:0];
  _RAND_2544 = {1{`RANDOM}};
  lineBuffer_2537 = _RAND_2544[7:0];
  _RAND_2545 = {1{`RANDOM}};
  lineBuffer_2538 = _RAND_2545[7:0];
  _RAND_2546 = {1{`RANDOM}};
  lineBuffer_2539 = _RAND_2546[7:0];
  _RAND_2547 = {1{`RANDOM}};
  lineBuffer_2540 = _RAND_2547[7:0];
  _RAND_2548 = {1{`RANDOM}};
  lineBuffer_2541 = _RAND_2548[7:0];
  _RAND_2549 = {1{`RANDOM}};
  lineBuffer_2542 = _RAND_2549[7:0];
  _RAND_2550 = {1{`RANDOM}};
  lineBuffer_2543 = _RAND_2550[7:0];
  _RAND_2551 = {1{`RANDOM}};
  lineBuffer_2544 = _RAND_2551[7:0];
  _RAND_2552 = {1{`RANDOM}};
  lineBuffer_2545 = _RAND_2552[7:0];
  _RAND_2553 = {1{`RANDOM}};
  lineBuffer_2546 = _RAND_2553[7:0];
  _RAND_2554 = {1{`RANDOM}};
  lineBuffer_2547 = _RAND_2554[7:0];
  _RAND_2555 = {1{`RANDOM}};
  lineBuffer_2548 = _RAND_2555[7:0];
  _RAND_2556 = {1{`RANDOM}};
  lineBuffer_2549 = _RAND_2556[7:0];
  _RAND_2557 = {1{`RANDOM}};
  lineBuffer_2550 = _RAND_2557[7:0];
  _RAND_2558 = {1{`RANDOM}};
  lineBuffer_2551 = _RAND_2558[7:0];
  _RAND_2559 = {1{`RANDOM}};
  lineBuffer_2552 = _RAND_2559[7:0];
  _RAND_2560 = {1{`RANDOM}};
  lineBuffer_2553 = _RAND_2560[7:0];
  _RAND_2561 = {1{`RANDOM}};
  lineBuffer_2554 = _RAND_2561[7:0];
  _RAND_2562 = {1{`RANDOM}};
  lineBuffer_2555 = _RAND_2562[7:0];
  _RAND_2563 = {1{`RANDOM}};
  lineBuffer_2556 = _RAND_2563[7:0];
  _RAND_2564 = {1{`RANDOM}};
  lineBuffer_2557 = _RAND_2564[7:0];
  _RAND_2565 = {1{`RANDOM}};
  lineBuffer_2558 = _RAND_2565[7:0];
  _RAND_2566 = {1{`RANDOM}};
  lineBuffer_2559 = _RAND_2566[7:0];
  _RAND_2567 = {1{`RANDOM}};
  lineBuffer_2560 = _RAND_2567[7:0];
  _RAND_2568 = {1{`RANDOM}};
  lineBuffer_2561 = _RAND_2568[7:0];
  _RAND_2569 = {1{`RANDOM}};
  lineBuffer_2562 = _RAND_2569[7:0];
  _RAND_2570 = {1{`RANDOM}};
  lineBuffer_2563 = _RAND_2570[7:0];
  _RAND_2571 = {1{`RANDOM}};
  lineBuffer_2564 = _RAND_2571[7:0];
  _RAND_2572 = {1{`RANDOM}};
  lineBuffer_2565 = _RAND_2572[7:0];
  _RAND_2573 = {1{`RANDOM}};
  lineBuffer_2566 = _RAND_2573[7:0];
  _RAND_2574 = {1{`RANDOM}};
  lineBuffer_2567 = _RAND_2574[7:0];
  _RAND_2575 = {1{`RANDOM}};
  lineBuffer_2568 = _RAND_2575[7:0];
  _RAND_2576 = {1{`RANDOM}};
  lineBuffer_2569 = _RAND_2576[7:0];
  _RAND_2577 = {1{`RANDOM}};
  lineBuffer_2570 = _RAND_2577[7:0];
  _RAND_2578 = {1{`RANDOM}};
  lineBuffer_2571 = _RAND_2578[7:0];
  _RAND_2579 = {1{`RANDOM}};
  lineBuffer_2572 = _RAND_2579[7:0];
  _RAND_2580 = {1{`RANDOM}};
  lineBuffer_2573 = _RAND_2580[7:0];
  _RAND_2581 = {1{`RANDOM}};
  lineBuffer_2574 = _RAND_2581[7:0];
  _RAND_2582 = {1{`RANDOM}};
  lineBuffer_2575 = _RAND_2582[7:0];
  _RAND_2583 = {1{`RANDOM}};
  lineBuffer_2576 = _RAND_2583[7:0];
  _RAND_2584 = {1{`RANDOM}};
  lineBuffer_2577 = _RAND_2584[7:0];
  _RAND_2585 = {1{`RANDOM}};
  lineBuffer_2578 = _RAND_2585[7:0];
  _RAND_2586 = {1{`RANDOM}};
  lineBuffer_2579 = _RAND_2586[7:0];
  _RAND_2587 = {1{`RANDOM}};
  lineBuffer_2580 = _RAND_2587[7:0];
  _RAND_2588 = {1{`RANDOM}};
  lineBuffer_2581 = _RAND_2588[7:0];
  _RAND_2589 = {1{`RANDOM}};
  lineBuffer_2582 = _RAND_2589[7:0];
  _RAND_2590 = {1{`RANDOM}};
  lineBuffer_2583 = _RAND_2590[7:0];
  _RAND_2591 = {1{`RANDOM}};
  lineBuffer_2584 = _RAND_2591[7:0];
  _RAND_2592 = {1{`RANDOM}};
  lineBuffer_2585 = _RAND_2592[7:0];
  _RAND_2593 = {1{`RANDOM}};
  lineBuffer_2586 = _RAND_2593[7:0];
  _RAND_2594 = {1{`RANDOM}};
  lineBuffer_2587 = _RAND_2594[7:0];
  _RAND_2595 = {1{`RANDOM}};
  lineBuffer_2588 = _RAND_2595[7:0];
  _RAND_2596 = {1{`RANDOM}};
  lineBuffer_2589 = _RAND_2596[7:0];
  _RAND_2597 = {1{`RANDOM}};
  lineBuffer_2590 = _RAND_2597[7:0];
  _RAND_2598 = {1{`RANDOM}};
  lineBuffer_2591 = _RAND_2598[7:0];
  _RAND_2599 = {1{`RANDOM}};
  lineBuffer_2592 = _RAND_2599[7:0];
  _RAND_2600 = {1{`RANDOM}};
  lineBuffer_2593 = _RAND_2600[7:0];
  _RAND_2601 = {1{`RANDOM}};
  lineBuffer_2594 = _RAND_2601[7:0];
  _RAND_2602 = {1{`RANDOM}};
  lineBuffer_2595 = _RAND_2602[7:0];
  _RAND_2603 = {1{`RANDOM}};
  lineBuffer_2596 = _RAND_2603[7:0];
  _RAND_2604 = {1{`RANDOM}};
  lineBuffer_2597 = _RAND_2604[7:0];
  _RAND_2605 = {1{`RANDOM}};
  lineBuffer_2598 = _RAND_2605[7:0];
  _RAND_2606 = {1{`RANDOM}};
  lineBuffer_2599 = _RAND_2606[7:0];
  _RAND_2607 = {1{`RANDOM}};
  lineBuffer_2600 = _RAND_2607[7:0];
  _RAND_2608 = {1{`RANDOM}};
  lineBuffer_2601 = _RAND_2608[7:0];
  _RAND_2609 = {1{`RANDOM}};
  lineBuffer_2602 = _RAND_2609[7:0];
  _RAND_2610 = {1{`RANDOM}};
  lineBuffer_2603 = _RAND_2610[7:0];
  _RAND_2611 = {1{`RANDOM}};
  lineBuffer_2604 = _RAND_2611[7:0];
  _RAND_2612 = {1{`RANDOM}};
  lineBuffer_2605 = _RAND_2612[7:0];
  _RAND_2613 = {1{`RANDOM}};
  lineBuffer_2606 = _RAND_2613[7:0];
  _RAND_2614 = {1{`RANDOM}};
  lineBuffer_2607 = _RAND_2614[7:0];
  _RAND_2615 = {1{`RANDOM}};
  lineBuffer_2608 = _RAND_2615[7:0];
  _RAND_2616 = {1{`RANDOM}};
  lineBuffer_2609 = _RAND_2616[7:0];
  _RAND_2617 = {1{`RANDOM}};
  lineBuffer_2610 = _RAND_2617[7:0];
  _RAND_2618 = {1{`RANDOM}};
  lineBuffer_2611 = _RAND_2618[7:0];
  _RAND_2619 = {1{`RANDOM}};
  lineBuffer_2612 = _RAND_2619[7:0];
  _RAND_2620 = {1{`RANDOM}};
  lineBuffer_2613 = _RAND_2620[7:0];
  _RAND_2621 = {1{`RANDOM}};
  lineBuffer_2614 = _RAND_2621[7:0];
  _RAND_2622 = {1{`RANDOM}};
  lineBuffer_2615 = _RAND_2622[7:0];
  _RAND_2623 = {1{`RANDOM}};
  lineBuffer_2616 = _RAND_2623[7:0];
  _RAND_2624 = {1{`RANDOM}};
  lineBuffer_2617 = _RAND_2624[7:0];
  _RAND_2625 = {1{`RANDOM}};
  lineBuffer_2618 = _RAND_2625[7:0];
  _RAND_2626 = {1{`RANDOM}};
  lineBuffer_2619 = _RAND_2626[7:0];
  _RAND_2627 = {1{`RANDOM}};
  lineBuffer_2620 = _RAND_2627[7:0];
  _RAND_2628 = {1{`RANDOM}};
  lineBuffer_2621 = _RAND_2628[7:0];
  _RAND_2629 = {1{`RANDOM}};
  lineBuffer_2622 = _RAND_2629[7:0];
  _RAND_2630 = {1{`RANDOM}};
  lineBuffer_2623 = _RAND_2630[7:0];
  _RAND_2631 = {1{`RANDOM}};
  lineBuffer_2624 = _RAND_2631[7:0];
  _RAND_2632 = {1{`RANDOM}};
  lineBuffer_2625 = _RAND_2632[7:0];
  _RAND_2633 = {1{`RANDOM}};
  lineBuffer_2626 = _RAND_2633[7:0];
  _RAND_2634 = {1{`RANDOM}};
  lineBuffer_2627 = _RAND_2634[7:0];
  _RAND_2635 = {1{`RANDOM}};
  lineBuffer_2628 = _RAND_2635[7:0];
  _RAND_2636 = {1{`RANDOM}};
  lineBuffer_2629 = _RAND_2636[7:0];
  _RAND_2637 = {1{`RANDOM}};
  lineBuffer_2630 = _RAND_2637[7:0];
  _RAND_2638 = {1{`RANDOM}};
  lineBuffer_2631 = _RAND_2638[7:0];
  _RAND_2639 = {1{`RANDOM}};
  lineBuffer_2632 = _RAND_2639[7:0];
  _RAND_2640 = {1{`RANDOM}};
  lineBuffer_2633 = _RAND_2640[7:0];
  _RAND_2641 = {1{`RANDOM}};
  lineBuffer_2634 = _RAND_2641[7:0];
  _RAND_2642 = {1{`RANDOM}};
  lineBuffer_2635 = _RAND_2642[7:0];
  _RAND_2643 = {1{`RANDOM}};
  lineBuffer_2636 = _RAND_2643[7:0];
  _RAND_2644 = {1{`RANDOM}};
  lineBuffer_2637 = _RAND_2644[7:0];
  _RAND_2645 = {1{`RANDOM}};
  lineBuffer_2638 = _RAND_2645[7:0];
  _RAND_2646 = {1{`RANDOM}};
  lineBuffer_2639 = _RAND_2646[7:0];
  _RAND_2647 = {1{`RANDOM}};
  lineBuffer_2640 = _RAND_2647[7:0];
  _RAND_2648 = {1{`RANDOM}};
  lineBuffer_2641 = _RAND_2648[7:0];
  _RAND_2649 = {1{`RANDOM}};
  lineBuffer_2642 = _RAND_2649[7:0];
  _RAND_2650 = {1{`RANDOM}};
  lineBuffer_2643 = _RAND_2650[7:0];
  _RAND_2651 = {1{`RANDOM}};
  lineBuffer_2644 = _RAND_2651[7:0];
  _RAND_2652 = {1{`RANDOM}};
  lineBuffer_2645 = _RAND_2652[7:0];
  _RAND_2653 = {1{`RANDOM}};
  lineBuffer_2646 = _RAND_2653[7:0];
  _RAND_2654 = {1{`RANDOM}};
  lineBuffer_2647 = _RAND_2654[7:0];
  _RAND_2655 = {1{`RANDOM}};
  lineBuffer_2648 = _RAND_2655[7:0];
  _RAND_2656 = {1{`RANDOM}};
  lineBuffer_2649 = _RAND_2656[7:0];
  _RAND_2657 = {1{`RANDOM}};
  lineBuffer_2650 = _RAND_2657[7:0];
  _RAND_2658 = {1{`RANDOM}};
  lineBuffer_2651 = _RAND_2658[7:0];
  _RAND_2659 = {1{`RANDOM}};
  lineBuffer_2652 = _RAND_2659[7:0];
  _RAND_2660 = {1{`RANDOM}};
  lineBuffer_2653 = _RAND_2660[7:0];
  _RAND_2661 = {1{`RANDOM}};
  lineBuffer_2654 = _RAND_2661[7:0];
  _RAND_2662 = {1{`RANDOM}};
  lineBuffer_2655 = _RAND_2662[7:0];
  _RAND_2663 = {1{`RANDOM}};
  lineBuffer_2656 = _RAND_2663[7:0];
  _RAND_2664 = {1{`RANDOM}};
  lineBuffer_2657 = _RAND_2664[7:0];
  _RAND_2665 = {1{`RANDOM}};
  lineBuffer_2658 = _RAND_2665[7:0];
  _RAND_2666 = {1{`RANDOM}};
  lineBuffer_2659 = _RAND_2666[7:0];
  _RAND_2667 = {1{`RANDOM}};
  lineBuffer_2660 = _RAND_2667[7:0];
  _RAND_2668 = {1{`RANDOM}};
  lineBuffer_2661 = _RAND_2668[7:0];
  _RAND_2669 = {1{`RANDOM}};
  lineBuffer_2662 = _RAND_2669[7:0];
  _RAND_2670 = {1{`RANDOM}};
  lineBuffer_2663 = _RAND_2670[7:0];
  _RAND_2671 = {1{`RANDOM}};
  lineBuffer_2664 = _RAND_2671[7:0];
  _RAND_2672 = {1{`RANDOM}};
  lineBuffer_2665 = _RAND_2672[7:0];
  _RAND_2673 = {1{`RANDOM}};
  lineBuffer_2666 = _RAND_2673[7:0];
  _RAND_2674 = {1{`RANDOM}};
  lineBuffer_2667 = _RAND_2674[7:0];
  _RAND_2675 = {1{`RANDOM}};
  lineBuffer_2668 = _RAND_2675[7:0];
  _RAND_2676 = {1{`RANDOM}};
  lineBuffer_2669 = _RAND_2676[7:0];
  _RAND_2677 = {1{`RANDOM}};
  lineBuffer_2670 = _RAND_2677[7:0];
  _RAND_2678 = {1{`RANDOM}};
  lineBuffer_2671 = _RAND_2678[7:0];
  _RAND_2679 = {1{`RANDOM}};
  lineBuffer_2672 = _RAND_2679[7:0];
  _RAND_2680 = {1{`RANDOM}};
  lineBuffer_2673 = _RAND_2680[7:0];
  _RAND_2681 = {1{`RANDOM}};
  lineBuffer_2674 = _RAND_2681[7:0];
  _RAND_2682 = {1{`RANDOM}};
  lineBuffer_2675 = _RAND_2682[7:0];
  _RAND_2683 = {1{`RANDOM}};
  lineBuffer_2676 = _RAND_2683[7:0];
  _RAND_2684 = {1{`RANDOM}};
  lineBuffer_2677 = _RAND_2684[7:0];
  _RAND_2685 = {1{`RANDOM}};
  lineBuffer_2678 = _RAND_2685[7:0];
  _RAND_2686 = {1{`RANDOM}};
  lineBuffer_2679 = _RAND_2686[7:0];
  _RAND_2687 = {1{`RANDOM}};
  lineBuffer_2680 = _RAND_2687[7:0];
  _RAND_2688 = {1{`RANDOM}};
  lineBuffer_2681 = _RAND_2688[7:0];
  _RAND_2689 = {1{`RANDOM}};
  lineBuffer_2682 = _RAND_2689[7:0];
  _RAND_2690 = {1{`RANDOM}};
  lineBuffer_2683 = _RAND_2690[7:0];
  _RAND_2691 = {1{`RANDOM}};
  lineBuffer_2684 = _RAND_2691[7:0];
  _RAND_2692 = {1{`RANDOM}};
  lineBuffer_2685 = _RAND_2692[7:0];
  _RAND_2693 = {1{`RANDOM}};
  lineBuffer_2686 = _RAND_2693[7:0];
  _RAND_2694 = {1{`RANDOM}};
  lineBuffer_2687 = _RAND_2694[7:0];
  _RAND_2695 = {1{`RANDOM}};
  lineBuffer_2688 = _RAND_2695[7:0];
  _RAND_2696 = {1{`RANDOM}};
  lineBuffer_2689 = _RAND_2696[7:0];
  _RAND_2697 = {1{`RANDOM}};
  lineBuffer_2690 = _RAND_2697[7:0];
  _RAND_2698 = {1{`RANDOM}};
  lineBuffer_2691 = _RAND_2698[7:0];
  _RAND_2699 = {1{`RANDOM}};
  lineBuffer_2692 = _RAND_2699[7:0];
  _RAND_2700 = {1{`RANDOM}};
  lineBuffer_2693 = _RAND_2700[7:0];
  _RAND_2701 = {1{`RANDOM}};
  lineBuffer_2694 = _RAND_2701[7:0];
  _RAND_2702 = {1{`RANDOM}};
  lineBuffer_2695 = _RAND_2702[7:0];
  _RAND_2703 = {1{`RANDOM}};
  lineBuffer_2696 = _RAND_2703[7:0];
  _RAND_2704 = {1{`RANDOM}};
  lineBuffer_2697 = _RAND_2704[7:0];
  _RAND_2705 = {1{`RANDOM}};
  lineBuffer_2698 = _RAND_2705[7:0];
  _RAND_2706 = {1{`RANDOM}};
  lineBuffer_2699 = _RAND_2706[7:0];
  _RAND_2707 = {1{`RANDOM}};
  lineBuffer_2700 = _RAND_2707[7:0];
  _RAND_2708 = {1{`RANDOM}};
  lineBuffer_2701 = _RAND_2708[7:0];
  _RAND_2709 = {1{`RANDOM}};
  lineBuffer_2702 = _RAND_2709[7:0];
  _RAND_2710 = {1{`RANDOM}};
  lineBuffer_2703 = _RAND_2710[7:0];
  _RAND_2711 = {1{`RANDOM}};
  lineBuffer_2704 = _RAND_2711[7:0];
  _RAND_2712 = {1{`RANDOM}};
  lineBuffer_2705 = _RAND_2712[7:0];
  _RAND_2713 = {1{`RANDOM}};
  lineBuffer_2706 = _RAND_2713[7:0];
  _RAND_2714 = {1{`RANDOM}};
  lineBuffer_2707 = _RAND_2714[7:0];
  _RAND_2715 = {1{`RANDOM}};
  lineBuffer_2708 = _RAND_2715[7:0];
  _RAND_2716 = {1{`RANDOM}};
  lineBuffer_2709 = _RAND_2716[7:0];
  _RAND_2717 = {1{`RANDOM}};
  lineBuffer_2710 = _RAND_2717[7:0];
  _RAND_2718 = {1{`RANDOM}};
  lineBuffer_2711 = _RAND_2718[7:0];
  _RAND_2719 = {1{`RANDOM}};
  lineBuffer_2712 = _RAND_2719[7:0];
  _RAND_2720 = {1{`RANDOM}};
  lineBuffer_2713 = _RAND_2720[7:0];
  _RAND_2721 = {1{`RANDOM}};
  lineBuffer_2714 = _RAND_2721[7:0];
  _RAND_2722 = {1{`RANDOM}};
  lineBuffer_2715 = _RAND_2722[7:0];
  _RAND_2723 = {1{`RANDOM}};
  lineBuffer_2716 = _RAND_2723[7:0];
  _RAND_2724 = {1{`RANDOM}};
  lineBuffer_2717 = _RAND_2724[7:0];
  _RAND_2725 = {1{`RANDOM}};
  lineBuffer_2718 = _RAND_2725[7:0];
  _RAND_2726 = {1{`RANDOM}};
  lineBuffer_2719 = _RAND_2726[7:0];
  _RAND_2727 = {1{`RANDOM}};
  lineBuffer_2720 = _RAND_2727[7:0];
  _RAND_2728 = {1{`RANDOM}};
  lineBuffer_2721 = _RAND_2728[7:0];
  _RAND_2729 = {1{`RANDOM}};
  lineBuffer_2722 = _RAND_2729[7:0];
  _RAND_2730 = {1{`RANDOM}};
  lineBuffer_2723 = _RAND_2730[7:0];
  _RAND_2731 = {1{`RANDOM}};
  lineBuffer_2724 = _RAND_2731[7:0];
  _RAND_2732 = {1{`RANDOM}};
  lineBuffer_2725 = _RAND_2732[7:0];
  _RAND_2733 = {1{`RANDOM}};
  lineBuffer_2726 = _RAND_2733[7:0];
  _RAND_2734 = {1{`RANDOM}};
  lineBuffer_2727 = _RAND_2734[7:0];
  _RAND_2735 = {1{`RANDOM}};
  lineBuffer_2728 = _RAND_2735[7:0];
  _RAND_2736 = {1{`RANDOM}};
  lineBuffer_2729 = _RAND_2736[7:0];
  _RAND_2737 = {1{`RANDOM}};
  lineBuffer_2730 = _RAND_2737[7:0];
  _RAND_2738 = {1{`RANDOM}};
  lineBuffer_2731 = _RAND_2738[7:0];
  _RAND_2739 = {1{`RANDOM}};
  lineBuffer_2732 = _RAND_2739[7:0];
  _RAND_2740 = {1{`RANDOM}};
  lineBuffer_2733 = _RAND_2740[7:0];
  _RAND_2741 = {1{`RANDOM}};
  lineBuffer_2734 = _RAND_2741[7:0];
  _RAND_2742 = {1{`RANDOM}};
  lineBuffer_2735 = _RAND_2742[7:0];
  _RAND_2743 = {1{`RANDOM}};
  lineBuffer_2736 = _RAND_2743[7:0];
  _RAND_2744 = {1{`RANDOM}};
  lineBuffer_2737 = _RAND_2744[7:0];
  _RAND_2745 = {1{`RANDOM}};
  lineBuffer_2738 = _RAND_2745[7:0];
  _RAND_2746 = {1{`RANDOM}};
  lineBuffer_2739 = _RAND_2746[7:0];
  _RAND_2747 = {1{`RANDOM}};
  lineBuffer_2740 = _RAND_2747[7:0];
  _RAND_2748 = {1{`RANDOM}};
  lineBuffer_2741 = _RAND_2748[7:0];
  _RAND_2749 = {1{`RANDOM}};
  lineBuffer_2742 = _RAND_2749[7:0];
  _RAND_2750 = {1{`RANDOM}};
  lineBuffer_2743 = _RAND_2750[7:0];
  _RAND_2751 = {1{`RANDOM}};
  lineBuffer_2744 = _RAND_2751[7:0];
  _RAND_2752 = {1{`RANDOM}};
  lineBuffer_2745 = _RAND_2752[7:0];
  _RAND_2753 = {1{`RANDOM}};
  lineBuffer_2746 = _RAND_2753[7:0];
  _RAND_2754 = {1{`RANDOM}};
  lineBuffer_2747 = _RAND_2754[7:0];
  _RAND_2755 = {1{`RANDOM}};
  lineBuffer_2748 = _RAND_2755[7:0];
  _RAND_2756 = {1{`RANDOM}};
  lineBuffer_2749 = _RAND_2756[7:0];
  _RAND_2757 = {1{`RANDOM}};
  lineBuffer_2750 = _RAND_2757[7:0];
  _RAND_2758 = {1{`RANDOM}};
  lineBuffer_2751 = _RAND_2758[7:0];
  _RAND_2759 = {1{`RANDOM}};
  lineBuffer_2752 = _RAND_2759[7:0];
  _RAND_2760 = {1{`RANDOM}};
  lineBuffer_2753 = _RAND_2760[7:0];
  _RAND_2761 = {1{`RANDOM}};
  lineBuffer_2754 = _RAND_2761[7:0];
  _RAND_2762 = {1{`RANDOM}};
  lineBuffer_2755 = _RAND_2762[7:0];
  _RAND_2763 = {1{`RANDOM}};
  lineBuffer_2756 = _RAND_2763[7:0];
  _RAND_2764 = {1{`RANDOM}};
  lineBuffer_2757 = _RAND_2764[7:0];
  _RAND_2765 = {1{`RANDOM}};
  lineBuffer_2758 = _RAND_2765[7:0];
  _RAND_2766 = {1{`RANDOM}};
  lineBuffer_2759 = _RAND_2766[7:0];
  _RAND_2767 = {1{`RANDOM}};
  lineBuffer_2760 = _RAND_2767[7:0];
  _RAND_2768 = {1{`RANDOM}};
  lineBuffer_2761 = _RAND_2768[7:0];
  _RAND_2769 = {1{`RANDOM}};
  lineBuffer_2762 = _RAND_2769[7:0];
  _RAND_2770 = {1{`RANDOM}};
  lineBuffer_2763 = _RAND_2770[7:0];
  _RAND_2771 = {1{`RANDOM}};
  lineBuffer_2764 = _RAND_2771[7:0];
  _RAND_2772 = {1{`RANDOM}};
  lineBuffer_2765 = _RAND_2772[7:0];
  _RAND_2773 = {1{`RANDOM}};
  lineBuffer_2766 = _RAND_2773[7:0];
  _RAND_2774 = {1{`RANDOM}};
  lineBuffer_2767 = _RAND_2774[7:0];
  _RAND_2775 = {1{`RANDOM}};
  lineBuffer_2768 = _RAND_2775[7:0];
  _RAND_2776 = {1{`RANDOM}};
  lineBuffer_2769 = _RAND_2776[7:0];
  _RAND_2777 = {1{`RANDOM}};
  lineBuffer_2770 = _RAND_2777[7:0];
  _RAND_2778 = {1{`RANDOM}};
  lineBuffer_2771 = _RAND_2778[7:0];
  _RAND_2779 = {1{`RANDOM}};
  lineBuffer_2772 = _RAND_2779[7:0];
  _RAND_2780 = {1{`RANDOM}};
  lineBuffer_2773 = _RAND_2780[7:0];
  _RAND_2781 = {1{`RANDOM}};
  lineBuffer_2774 = _RAND_2781[7:0];
  _RAND_2782 = {1{`RANDOM}};
  lineBuffer_2775 = _RAND_2782[7:0];
  _RAND_2783 = {1{`RANDOM}};
  lineBuffer_2776 = _RAND_2783[7:0];
  _RAND_2784 = {1{`RANDOM}};
  lineBuffer_2777 = _RAND_2784[7:0];
  _RAND_2785 = {1{`RANDOM}};
  lineBuffer_2778 = _RAND_2785[7:0];
  _RAND_2786 = {1{`RANDOM}};
  lineBuffer_2779 = _RAND_2786[7:0];
  _RAND_2787 = {1{`RANDOM}};
  lineBuffer_2780 = _RAND_2787[7:0];
  _RAND_2788 = {1{`RANDOM}};
  lineBuffer_2781 = _RAND_2788[7:0];
  _RAND_2789 = {1{`RANDOM}};
  lineBuffer_2782 = _RAND_2789[7:0];
  _RAND_2790 = {1{`RANDOM}};
  lineBuffer_2783 = _RAND_2790[7:0];
  _RAND_2791 = {1{`RANDOM}};
  lineBuffer_2784 = _RAND_2791[7:0];
  _RAND_2792 = {1{`RANDOM}};
  lineBuffer_2785 = _RAND_2792[7:0];
  _RAND_2793 = {1{`RANDOM}};
  lineBuffer_2786 = _RAND_2793[7:0];
  _RAND_2794 = {1{`RANDOM}};
  lineBuffer_2787 = _RAND_2794[7:0];
  _RAND_2795 = {1{`RANDOM}};
  lineBuffer_2788 = _RAND_2795[7:0];
  _RAND_2796 = {1{`RANDOM}};
  lineBuffer_2789 = _RAND_2796[7:0];
  _RAND_2797 = {1{`RANDOM}};
  lineBuffer_2790 = _RAND_2797[7:0];
  _RAND_2798 = {1{`RANDOM}};
  lineBuffer_2791 = _RAND_2798[7:0];
  _RAND_2799 = {1{`RANDOM}};
  lineBuffer_2792 = _RAND_2799[7:0];
  _RAND_2800 = {1{`RANDOM}};
  lineBuffer_2793 = _RAND_2800[7:0];
  _RAND_2801 = {1{`RANDOM}};
  lineBuffer_2794 = _RAND_2801[7:0];
  _RAND_2802 = {1{`RANDOM}};
  lineBuffer_2795 = _RAND_2802[7:0];
  _RAND_2803 = {1{`RANDOM}};
  lineBuffer_2796 = _RAND_2803[7:0];
  _RAND_2804 = {1{`RANDOM}};
  lineBuffer_2797 = _RAND_2804[7:0];
  _RAND_2805 = {1{`RANDOM}};
  lineBuffer_2798 = _RAND_2805[7:0];
  _RAND_2806 = {1{`RANDOM}};
  lineBuffer_2799 = _RAND_2806[7:0];
  _RAND_2807 = {1{`RANDOM}};
  lineBuffer_2800 = _RAND_2807[7:0];
  _RAND_2808 = {1{`RANDOM}};
  lineBuffer_2801 = _RAND_2808[7:0];
  _RAND_2809 = {1{`RANDOM}};
  lineBuffer_2802 = _RAND_2809[7:0];
  _RAND_2810 = {1{`RANDOM}};
  lineBuffer_2803 = _RAND_2810[7:0];
  _RAND_2811 = {1{`RANDOM}};
  lineBuffer_2804 = _RAND_2811[7:0];
  _RAND_2812 = {1{`RANDOM}};
  lineBuffer_2805 = _RAND_2812[7:0];
  _RAND_2813 = {1{`RANDOM}};
  lineBuffer_2806 = _RAND_2813[7:0];
  _RAND_2814 = {1{`RANDOM}};
  lineBuffer_2807 = _RAND_2814[7:0];
  _RAND_2815 = {1{`RANDOM}};
  lineBuffer_2808 = _RAND_2815[7:0];
  _RAND_2816 = {1{`RANDOM}};
  lineBuffer_2809 = _RAND_2816[7:0];
  _RAND_2817 = {1{`RANDOM}};
  lineBuffer_2810 = _RAND_2817[7:0];
  _RAND_2818 = {1{`RANDOM}};
  lineBuffer_2811 = _RAND_2818[7:0];
  _RAND_2819 = {1{`RANDOM}};
  lineBuffer_2812 = _RAND_2819[7:0];
  _RAND_2820 = {1{`RANDOM}};
  lineBuffer_2813 = _RAND_2820[7:0];
  _RAND_2821 = {1{`RANDOM}};
  lineBuffer_2814 = _RAND_2821[7:0];
  _RAND_2822 = {1{`RANDOM}};
  lineBuffer_2815 = _RAND_2822[7:0];
  _RAND_2823 = {1{`RANDOM}};
  lineBuffer_2816 = _RAND_2823[7:0];
  _RAND_2824 = {1{`RANDOM}};
  lineBuffer_2817 = _RAND_2824[7:0];
  _RAND_2825 = {1{`RANDOM}};
  lineBuffer_2818 = _RAND_2825[7:0];
  _RAND_2826 = {1{`RANDOM}};
  lineBuffer_2819 = _RAND_2826[7:0];
  _RAND_2827 = {1{`RANDOM}};
  lineBuffer_2820 = _RAND_2827[7:0];
  _RAND_2828 = {1{`RANDOM}};
  lineBuffer_2821 = _RAND_2828[7:0];
  _RAND_2829 = {1{`RANDOM}};
  lineBuffer_2822 = _RAND_2829[7:0];
  _RAND_2830 = {1{`RANDOM}};
  lineBuffer_2823 = _RAND_2830[7:0];
  _RAND_2831 = {1{`RANDOM}};
  lineBuffer_2824 = _RAND_2831[7:0];
  _RAND_2832 = {1{`RANDOM}};
  lineBuffer_2825 = _RAND_2832[7:0];
  _RAND_2833 = {1{`RANDOM}};
  lineBuffer_2826 = _RAND_2833[7:0];
  _RAND_2834 = {1{`RANDOM}};
  lineBuffer_2827 = _RAND_2834[7:0];
  _RAND_2835 = {1{`RANDOM}};
  lineBuffer_2828 = _RAND_2835[7:0];
  _RAND_2836 = {1{`RANDOM}};
  lineBuffer_2829 = _RAND_2836[7:0];
  _RAND_2837 = {1{`RANDOM}};
  lineBuffer_2830 = _RAND_2837[7:0];
  _RAND_2838 = {1{`RANDOM}};
  lineBuffer_2831 = _RAND_2838[7:0];
  _RAND_2839 = {1{`RANDOM}};
  lineBuffer_2832 = _RAND_2839[7:0];
  _RAND_2840 = {1{`RANDOM}};
  lineBuffer_2833 = _RAND_2840[7:0];
  _RAND_2841 = {1{`RANDOM}};
  lineBuffer_2834 = _RAND_2841[7:0];
  _RAND_2842 = {1{`RANDOM}};
  lineBuffer_2835 = _RAND_2842[7:0];
  _RAND_2843 = {1{`RANDOM}};
  lineBuffer_2836 = _RAND_2843[7:0];
  _RAND_2844 = {1{`RANDOM}};
  lineBuffer_2837 = _RAND_2844[7:0];
  _RAND_2845 = {1{`RANDOM}};
  lineBuffer_2838 = _RAND_2845[7:0];
  _RAND_2846 = {1{`RANDOM}};
  lineBuffer_2839 = _RAND_2846[7:0];
  _RAND_2847 = {1{`RANDOM}};
  lineBuffer_2840 = _RAND_2847[7:0];
  _RAND_2848 = {1{`RANDOM}};
  lineBuffer_2841 = _RAND_2848[7:0];
  _RAND_2849 = {1{`RANDOM}};
  lineBuffer_2842 = _RAND_2849[7:0];
  _RAND_2850 = {1{`RANDOM}};
  lineBuffer_2843 = _RAND_2850[7:0];
  _RAND_2851 = {1{`RANDOM}};
  lineBuffer_2844 = _RAND_2851[7:0];
  _RAND_2852 = {1{`RANDOM}};
  lineBuffer_2845 = _RAND_2852[7:0];
  _RAND_2853 = {1{`RANDOM}};
  lineBuffer_2846 = _RAND_2853[7:0];
  _RAND_2854 = {1{`RANDOM}};
  lineBuffer_2847 = _RAND_2854[7:0];
  _RAND_2855 = {1{`RANDOM}};
  lineBuffer_2848 = _RAND_2855[7:0];
  _RAND_2856 = {1{`RANDOM}};
  lineBuffer_2849 = _RAND_2856[7:0];
  _RAND_2857 = {1{`RANDOM}};
  lineBuffer_2850 = _RAND_2857[7:0];
  _RAND_2858 = {1{`RANDOM}};
  lineBuffer_2851 = _RAND_2858[7:0];
  _RAND_2859 = {1{`RANDOM}};
  lineBuffer_2852 = _RAND_2859[7:0];
  _RAND_2860 = {1{`RANDOM}};
  lineBuffer_2853 = _RAND_2860[7:0];
  _RAND_2861 = {1{`RANDOM}};
  lineBuffer_2854 = _RAND_2861[7:0];
  _RAND_2862 = {1{`RANDOM}};
  lineBuffer_2855 = _RAND_2862[7:0];
  _RAND_2863 = {1{`RANDOM}};
  lineBuffer_2856 = _RAND_2863[7:0];
  _RAND_2864 = {1{`RANDOM}};
  lineBuffer_2857 = _RAND_2864[7:0];
  _RAND_2865 = {1{`RANDOM}};
  lineBuffer_2858 = _RAND_2865[7:0];
  _RAND_2866 = {1{`RANDOM}};
  lineBuffer_2859 = _RAND_2866[7:0];
  _RAND_2867 = {1{`RANDOM}};
  lineBuffer_2860 = _RAND_2867[7:0];
  _RAND_2868 = {1{`RANDOM}};
  lineBuffer_2861 = _RAND_2868[7:0];
  _RAND_2869 = {1{`RANDOM}};
  lineBuffer_2862 = _RAND_2869[7:0];
  _RAND_2870 = {1{`RANDOM}};
  lineBuffer_2863 = _RAND_2870[7:0];
  _RAND_2871 = {1{`RANDOM}};
  lineBuffer_2864 = _RAND_2871[7:0];
  _RAND_2872 = {1{`RANDOM}};
  lineBuffer_2865 = _RAND_2872[7:0];
  _RAND_2873 = {1{`RANDOM}};
  lineBuffer_2866 = _RAND_2873[7:0];
  _RAND_2874 = {1{`RANDOM}};
  lineBuffer_2867 = _RAND_2874[7:0];
  _RAND_2875 = {1{`RANDOM}};
  lineBuffer_2868 = _RAND_2875[7:0];
  _RAND_2876 = {1{`RANDOM}};
  lineBuffer_2869 = _RAND_2876[7:0];
  _RAND_2877 = {1{`RANDOM}};
  lineBuffer_2870 = _RAND_2877[7:0];
  _RAND_2878 = {1{`RANDOM}};
  lineBuffer_2871 = _RAND_2878[7:0];
  _RAND_2879 = {1{`RANDOM}};
  lineBuffer_2872 = _RAND_2879[7:0];
  _RAND_2880 = {1{`RANDOM}};
  lineBuffer_2873 = _RAND_2880[7:0];
  _RAND_2881 = {1{`RANDOM}};
  lineBuffer_2874 = _RAND_2881[7:0];
  _RAND_2882 = {1{`RANDOM}};
  lineBuffer_2875 = _RAND_2882[7:0];
  _RAND_2883 = {1{`RANDOM}};
  lineBuffer_2876 = _RAND_2883[7:0];
  _RAND_2884 = {1{`RANDOM}};
  lineBuffer_2877 = _RAND_2884[7:0];
  _RAND_2885 = {1{`RANDOM}};
  lineBuffer_2878 = _RAND_2885[7:0];
  _RAND_2886 = {1{`RANDOM}};
  lineBuffer_2879 = _RAND_2886[7:0];
  _RAND_2887 = {1{`RANDOM}};
  lineBuffer_2880 = _RAND_2887[7:0];
  _RAND_2888 = {1{`RANDOM}};
  lineBuffer_2881 = _RAND_2888[7:0];
  _RAND_2889 = {1{`RANDOM}};
  lineBuffer_2882 = _RAND_2889[7:0];
  _RAND_2890 = {1{`RANDOM}};
  lineBuffer_2883 = _RAND_2890[7:0];
  _RAND_2891 = {1{`RANDOM}};
  lineBuffer_2884 = _RAND_2891[7:0];
  _RAND_2892 = {1{`RANDOM}};
  lineBuffer_2885 = _RAND_2892[7:0];
  _RAND_2893 = {1{`RANDOM}};
  lineBuffer_2886 = _RAND_2893[7:0];
  _RAND_2894 = {1{`RANDOM}};
  lineBuffer_2887 = _RAND_2894[7:0];
  _RAND_2895 = {1{`RANDOM}};
  lineBuffer_2888 = _RAND_2895[7:0];
  _RAND_2896 = {1{`RANDOM}};
  lineBuffer_2889 = _RAND_2896[7:0];
  _RAND_2897 = {1{`RANDOM}};
  lineBuffer_2890 = _RAND_2897[7:0];
  _RAND_2898 = {1{`RANDOM}};
  lineBuffer_2891 = _RAND_2898[7:0];
  _RAND_2899 = {1{`RANDOM}};
  lineBuffer_2892 = _RAND_2899[7:0];
  _RAND_2900 = {1{`RANDOM}};
  lineBuffer_2893 = _RAND_2900[7:0];
  _RAND_2901 = {1{`RANDOM}};
  lineBuffer_2894 = _RAND_2901[7:0];
  _RAND_2902 = {1{`RANDOM}};
  lineBuffer_2895 = _RAND_2902[7:0];
  _RAND_2903 = {1{`RANDOM}};
  lineBuffer_2896 = _RAND_2903[7:0];
  _RAND_2904 = {1{`RANDOM}};
  lineBuffer_2897 = _RAND_2904[7:0];
  _RAND_2905 = {1{`RANDOM}};
  lineBuffer_2898 = _RAND_2905[7:0];
  _RAND_2906 = {1{`RANDOM}};
  lineBuffer_2899 = _RAND_2906[7:0];
  _RAND_2907 = {1{`RANDOM}};
  lineBuffer_2900 = _RAND_2907[7:0];
  _RAND_2908 = {1{`RANDOM}};
  lineBuffer_2901 = _RAND_2908[7:0];
  _RAND_2909 = {1{`RANDOM}};
  lineBuffer_2902 = _RAND_2909[7:0];
  _RAND_2910 = {1{`RANDOM}};
  lineBuffer_2903 = _RAND_2910[7:0];
  _RAND_2911 = {1{`RANDOM}};
  lineBuffer_2904 = _RAND_2911[7:0];
  _RAND_2912 = {1{`RANDOM}};
  lineBuffer_2905 = _RAND_2912[7:0];
  _RAND_2913 = {1{`RANDOM}};
  lineBuffer_2906 = _RAND_2913[7:0];
  _RAND_2914 = {1{`RANDOM}};
  lineBuffer_2907 = _RAND_2914[7:0];
  _RAND_2915 = {1{`RANDOM}};
  lineBuffer_2908 = _RAND_2915[7:0];
  _RAND_2916 = {1{`RANDOM}};
  lineBuffer_2909 = _RAND_2916[7:0];
  _RAND_2917 = {1{`RANDOM}};
  lineBuffer_2910 = _RAND_2917[7:0];
  _RAND_2918 = {1{`RANDOM}};
  lineBuffer_2911 = _RAND_2918[7:0];
  _RAND_2919 = {1{`RANDOM}};
  lineBuffer_2912 = _RAND_2919[7:0];
  _RAND_2920 = {1{`RANDOM}};
  lineBuffer_2913 = _RAND_2920[7:0];
  _RAND_2921 = {1{`RANDOM}};
  lineBuffer_2914 = _RAND_2921[7:0];
  _RAND_2922 = {1{`RANDOM}};
  lineBuffer_2915 = _RAND_2922[7:0];
  _RAND_2923 = {1{`RANDOM}};
  lineBuffer_2916 = _RAND_2923[7:0];
  _RAND_2924 = {1{`RANDOM}};
  lineBuffer_2917 = _RAND_2924[7:0];
  _RAND_2925 = {1{`RANDOM}};
  lineBuffer_2918 = _RAND_2925[7:0];
  _RAND_2926 = {1{`RANDOM}};
  lineBuffer_2919 = _RAND_2926[7:0];
  _RAND_2927 = {1{`RANDOM}};
  lineBuffer_2920 = _RAND_2927[7:0];
  _RAND_2928 = {1{`RANDOM}};
  lineBuffer_2921 = _RAND_2928[7:0];
  _RAND_2929 = {1{`RANDOM}};
  lineBuffer_2922 = _RAND_2929[7:0];
  _RAND_2930 = {1{`RANDOM}};
  lineBuffer_2923 = _RAND_2930[7:0];
  _RAND_2931 = {1{`RANDOM}};
  lineBuffer_2924 = _RAND_2931[7:0];
  _RAND_2932 = {1{`RANDOM}};
  lineBuffer_2925 = _RAND_2932[7:0];
  _RAND_2933 = {1{`RANDOM}};
  lineBuffer_2926 = _RAND_2933[7:0];
  _RAND_2934 = {1{`RANDOM}};
  lineBuffer_2927 = _RAND_2934[7:0];
  _RAND_2935 = {1{`RANDOM}};
  lineBuffer_2928 = _RAND_2935[7:0];
  _RAND_2936 = {1{`RANDOM}};
  lineBuffer_2929 = _RAND_2936[7:0];
  _RAND_2937 = {1{`RANDOM}};
  lineBuffer_2930 = _RAND_2937[7:0];
  _RAND_2938 = {1{`RANDOM}};
  lineBuffer_2931 = _RAND_2938[7:0];
  _RAND_2939 = {1{`RANDOM}};
  lineBuffer_2932 = _RAND_2939[7:0];
  _RAND_2940 = {1{`RANDOM}};
  lineBuffer_2933 = _RAND_2940[7:0];
  _RAND_2941 = {1{`RANDOM}};
  lineBuffer_2934 = _RAND_2941[7:0];
  _RAND_2942 = {1{`RANDOM}};
  lineBuffer_2935 = _RAND_2942[7:0];
  _RAND_2943 = {1{`RANDOM}};
  lineBuffer_2936 = _RAND_2943[7:0];
  _RAND_2944 = {1{`RANDOM}};
  lineBuffer_2937 = _RAND_2944[7:0];
  _RAND_2945 = {1{`RANDOM}};
  lineBuffer_2938 = _RAND_2945[7:0];
  _RAND_2946 = {1{`RANDOM}};
  lineBuffer_2939 = _RAND_2946[7:0];
  _RAND_2947 = {1{`RANDOM}};
  lineBuffer_2940 = _RAND_2947[7:0];
  _RAND_2948 = {1{`RANDOM}};
  lineBuffer_2941 = _RAND_2948[7:0];
  _RAND_2949 = {1{`RANDOM}};
  lineBuffer_2942 = _RAND_2949[7:0];
  _RAND_2950 = {1{`RANDOM}};
  lineBuffer_2943 = _RAND_2950[7:0];
  _RAND_2951 = {1{`RANDOM}};
  lineBuffer_2944 = _RAND_2951[7:0];
  _RAND_2952 = {1{`RANDOM}};
  lineBuffer_2945 = _RAND_2952[7:0];
  _RAND_2953 = {1{`RANDOM}};
  lineBuffer_2946 = _RAND_2953[7:0];
  _RAND_2954 = {1{`RANDOM}};
  lineBuffer_2947 = _RAND_2954[7:0];
  _RAND_2955 = {1{`RANDOM}};
  lineBuffer_2948 = _RAND_2955[7:0];
  _RAND_2956 = {1{`RANDOM}};
  lineBuffer_2949 = _RAND_2956[7:0];
  _RAND_2957 = {1{`RANDOM}};
  lineBuffer_2950 = _RAND_2957[7:0];
  _RAND_2958 = {1{`RANDOM}};
  lineBuffer_2951 = _RAND_2958[7:0];
  _RAND_2959 = {1{`RANDOM}};
  lineBuffer_2952 = _RAND_2959[7:0];
  _RAND_2960 = {1{`RANDOM}};
  lineBuffer_2953 = _RAND_2960[7:0];
  _RAND_2961 = {1{`RANDOM}};
  lineBuffer_2954 = _RAND_2961[7:0];
  _RAND_2962 = {1{`RANDOM}};
  lineBuffer_2955 = _RAND_2962[7:0];
  _RAND_2963 = {1{`RANDOM}};
  lineBuffer_2956 = _RAND_2963[7:0];
  _RAND_2964 = {1{`RANDOM}};
  lineBuffer_2957 = _RAND_2964[7:0];
  _RAND_2965 = {1{`RANDOM}};
  lineBuffer_2958 = _RAND_2965[7:0];
  _RAND_2966 = {1{`RANDOM}};
  lineBuffer_2959 = _RAND_2966[7:0];
  _RAND_2967 = {1{`RANDOM}};
  lineBuffer_2960 = _RAND_2967[7:0];
  _RAND_2968 = {1{`RANDOM}};
  lineBuffer_2961 = _RAND_2968[7:0];
  _RAND_2969 = {1{`RANDOM}};
  lineBuffer_2962 = _RAND_2969[7:0];
  _RAND_2970 = {1{`RANDOM}};
  lineBuffer_2963 = _RAND_2970[7:0];
  _RAND_2971 = {1{`RANDOM}};
  lineBuffer_2964 = _RAND_2971[7:0];
  _RAND_2972 = {1{`RANDOM}};
  lineBuffer_2965 = _RAND_2972[7:0];
  _RAND_2973 = {1{`RANDOM}};
  lineBuffer_2966 = _RAND_2973[7:0];
  _RAND_2974 = {1{`RANDOM}};
  lineBuffer_2967 = _RAND_2974[7:0];
  _RAND_2975 = {1{`RANDOM}};
  lineBuffer_2968 = _RAND_2975[7:0];
  _RAND_2976 = {1{`RANDOM}};
  lineBuffer_2969 = _RAND_2976[7:0];
  _RAND_2977 = {1{`RANDOM}};
  lineBuffer_2970 = _RAND_2977[7:0];
  _RAND_2978 = {1{`RANDOM}};
  lineBuffer_2971 = _RAND_2978[7:0];
  _RAND_2979 = {1{`RANDOM}};
  lineBuffer_2972 = _RAND_2979[7:0];
  _RAND_2980 = {1{`RANDOM}};
  lineBuffer_2973 = _RAND_2980[7:0];
  _RAND_2981 = {1{`RANDOM}};
  lineBuffer_2974 = _RAND_2981[7:0];
  _RAND_2982 = {1{`RANDOM}};
  lineBuffer_2975 = _RAND_2982[7:0];
  _RAND_2983 = {1{`RANDOM}};
  lineBuffer_2976 = _RAND_2983[7:0];
  _RAND_2984 = {1{`RANDOM}};
  lineBuffer_2977 = _RAND_2984[7:0];
  _RAND_2985 = {1{`RANDOM}};
  lineBuffer_2978 = _RAND_2985[7:0];
  _RAND_2986 = {1{`RANDOM}};
  lineBuffer_2979 = _RAND_2986[7:0];
  _RAND_2987 = {1{`RANDOM}};
  lineBuffer_2980 = _RAND_2987[7:0];
  _RAND_2988 = {1{`RANDOM}};
  lineBuffer_2981 = _RAND_2988[7:0];
  _RAND_2989 = {1{`RANDOM}};
  lineBuffer_2982 = _RAND_2989[7:0];
  _RAND_2990 = {1{`RANDOM}};
  lineBuffer_2983 = _RAND_2990[7:0];
  _RAND_2991 = {1{`RANDOM}};
  lineBuffer_2984 = _RAND_2991[7:0];
  _RAND_2992 = {1{`RANDOM}};
  lineBuffer_2985 = _RAND_2992[7:0];
  _RAND_2993 = {1{`RANDOM}};
  lineBuffer_2986 = _RAND_2993[7:0];
  _RAND_2994 = {1{`RANDOM}};
  lineBuffer_2987 = _RAND_2994[7:0];
  _RAND_2995 = {1{`RANDOM}};
  lineBuffer_2988 = _RAND_2995[7:0];
  _RAND_2996 = {1{`RANDOM}};
  lineBuffer_2989 = _RAND_2996[7:0];
  _RAND_2997 = {1{`RANDOM}};
  lineBuffer_2990 = _RAND_2997[7:0];
  _RAND_2998 = {1{`RANDOM}};
  lineBuffer_2991 = _RAND_2998[7:0];
  _RAND_2999 = {1{`RANDOM}};
  lineBuffer_2992 = _RAND_2999[7:0];
  _RAND_3000 = {1{`RANDOM}};
  lineBuffer_2993 = _RAND_3000[7:0];
  _RAND_3001 = {1{`RANDOM}};
  lineBuffer_2994 = _RAND_3001[7:0];
  _RAND_3002 = {1{`RANDOM}};
  lineBuffer_2995 = _RAND_3002[7:0];
  _RAND_3003 = {1{`RANDOM}};
  lineBuffer_2996 = _RAND_3003[7:0];
  _RAND_3004 = {1{`RANDOM}};
  lineBuffer_2997 = _RAND_3004[7:0];
  _RAND_3005 = {1{`RANDOM}};
  lineBuffer_2998 = _RAND_3005[7:0];
  _RAND_3006 = {1{`RANDOM}};
  lineBuffer_2999 = _RAND_3006[7:0];
  _RAND_3007 = {1{`RANDOM}};
  lineBuffer_3000 = _RAND_3007[7:0];
  _RAND_3008 = {1{`RANDOM}};
  lineBuffer_3001 = _RAND_3008[7:0];
  _RAND_3009 = {1{`RANDOM}};
  lineBuffer_3002 = _RAND_3009[7:0];
  _RAND_3010 = {1{`RANDOM}};
  lineBuffer_3003 = _RAND_3010[7:0];
  _RAND_3011 = {1{`RANDOM}};
  lineBuffer_3004 = _RAND_3011[7:0];
  _RAND_3012 = {1{`RANDOM}};
  lineBuffer_3005 = _RAND_3012[7:0];
  _RAND_3013 = {1{`RANDOM}};
  lineBuffer_3006 = _RAND_3013[7:0];
  _RAND_3014 = {1{`RANDOM}};
  lineBuffer_3007 = _RAND_3014[7:0];
  _RAND_3015 = {1{`RANDOM}};
  lineBuffer_3008 = _RAND_3015[7:0];
  _RAND_3016 = {1{`RANDOM}};
  lineBuffer_3009 = _RAND_3016[7:0];
  _RAND_3017 = {1{`RANDOM}};
  lineBuffer_3010 = _RAND_3017[7:0];
  _RAND_3018 = {1{`RANDOM}};
  lineBuffer_3011 = _RAND_3018[7:0];
  _RAND_3019 = {1{`RANDOM}};
  lineBuffer_3012 = _RAND_3019[7:0];
  _RAND_3020 = {1{`RANDOM}};
  lineBuffer_3013 = _RAND_3020[7:0];
  _RAND_3021 = {1{`RANDOM}};
  lineBuffer_3014 = _RAND_3021[7:0];
  _RAND_3022 = {1{`RANDOM}};
  lineBuffer_3015 = _RAND_3022[7:0];
  _RAND_3023 = {1{`RANDOM}};
  lineBuffer_3016 = _RAND_3023[7:0];
  _RAND_3024 = {1{`RANDOM}};
  lineBuffer_3017 = _RAND_3024[7:0];
  _RAND_3025 = {1{`RANDOM}};
  lineBuffer_3018 = _RAND_3025[7:0];
  _RAND_3026 = {1{`RANDOM}};
  lineBuffer_3019 = _RAND_3026[7:0];
  _RAND_3027 = {1{`RANDOM}};
  lineBuffer_3020 = _RAND_3027[7:0];
  _RAND_3028 = {1{`RANDOM}};
  lineBuffer_3021 = _RAND_3028[7:0];
  _RAND_3029 = {1{`RANDOM}};
  lineBuffer_3022 = _RAND_3029[7:0];
  _RAND_3030 = {1{`RANDOM}};
  lineBuffer_3023 = _RAND_3030[7:0];
  _RAND_3031 = {1{`RANDOM}};
  lineBuffer_3024 = _RAND_3031[7:0];
  _RAND_3032 = {1{`RANDOM}};
  lineBuffer_3025 = _RAND_3032[7:0];
  _RAND_3033 = {1{`RANDOM}};
  lineBuffer_3026 = _RAND_3033[7:0];
  _RAND_3034 = {1{`RANDOM}};
  lineBuffer_3027 = _RAND_3034[7:0];
  _RAND_3035 = {1{`RANDOM}};
  lineBuffer_3028 = _RAND_3035[7:0];
  _RAND_3036 = {1{`RANDOM}};
  lineBuffer_3029 = _RAND_3036[7:0];
  _RAND_3037 = {1{`RANDOM}};
  lineBuffer_3030 = _RAND_3037[7:0];
  _RAND_3038 = {1{`RANDOM}};
  lineBuffer_3031 = _RAND_3038[7:0];
  _RAND_3039 = {1{`RANDOM}};
  lineBuffer_3032 = _RAND_3039[7:0];
  _RAND_3040 = {1{`RANDOM}};
  lineBuffer_3033 = _RAND_3040[7:0];
  _RAND_3041 = {1{`RANDOM}};
  lineBuffer_3034 = _RAND_3041[7:0];
  _RAND_3042 = {1{`RANDOM}};
  lineBuffer_3035 = _RAND_3042[7:0];
  _RAND_3043 = {1{`RANDOM}};
  lineBuffer_3036 = _RAND_3043[7:0];
  _RAND_3044 = {1{`RANDOM}};
  lineBuffer_3037 = _RAND_3044[7:0];
  _RAND_3045 = {1{`RANDOM}};
  lineBuffer_3038 = _RAND_3045[7:0];
  _RAND_3046 = {1{`RANDOM}};
  lineBuffer_3039 = _RAND_3046[7:0];
  _RAND_3047 = {1{`RANDOM}};
  lineBuffer_3040 = _RAND_3047[7:0];
  _RAND_3048 = {1{`RANDOM}};
  lineBuffer_3041 = _RAND_3048[7:0];
  _RAND_3049 = {1{`RANDOM}};
  lineBuffer_3042 = _RAND_3049[7:0];
  _RAND_3050 = {1{`RANDOM}};
  lineBuffer_3043 = _RAND_3050[7:0];
  _RAND_3051 = {1{`RANDOM}};
  lineBuffer_3044 = _RAND_3051[7:0];
  _RAND_3052 = {1{`RANDOM}};
  lineBuffer_3045 = _RAND_3052[7:0];
  _RAND_3053 = {1{`RANDOM}};
  lineBuffer_3046 = _RAND_3053[7:0];
  _RAND_3054 = {1{`RANDOM}};
  lineBuffer_3047 = _RAND_3054[7:0];
  _RAND_3055 = {1{`RANDOM}};
  lineBuffer_3048 = _RAND_3055[7:0];
  _RAND_3056 = {1{`RANDOM}};
  lineBuffer_3049 = _RAND_3056[7:0];
  _RAND_3057 = {1{`RANDOM}};
  lineBuffer_3050 = _RAND_3057[7:0];
  _RAND_3058 = {1{`RANDOM}};
  lineBuffer_3051 = _RAND_3058[7:0];
  _RAND_3059 = {1{`RANDOM}};
  lineBuffer_3052 = _RAND_3059[7:0];
  _RAND_3060 = {1{`RANDOM}};
  lineBuffer_3053 = _RAND_3060[7:0];
  _RAND_3061 = {1{`RANDOM}};
  lineBuffer_3054 = _RAND_3061[7:0];
  _RAND_3062 = {1{`RANDOM}};
  lineBuffer_3055 = _RAND_3062[7:0];
  _RAND_3063 = {1{`RANDOM}};
  lineBuffer_3056 = _RAND_3063[7:0];
  _RAND_3064 = {1{`RANDOM}};
  lineBuffer_3057 = _RAND_3064[7:0];
  _RAND_3065 = {1{`RANDOM}};
  lineBuffer_3058 = _RAND_3065[7:0];
  _RAND_3066 = {1{`RANDOM}};
  lineBuffer_3059 = _RAND_3066[7:0];
  _RAND_3067 = {1{`RANDOM}};
  lineBuffer_3060 = _RAND_3067[7:0];
  _RAND_3068 = {1{`RANDOM}};
  lineBuffer_3061 = _RAND_3068[7:0];
  _RAND_3069 = {1{`RANDOM}};
  lineBuffer_3062 = _RAND_3069[7:0];
  _RAND_3070 = {1{`RANDOM}};
  lineBuffer_3063 = _RAND_3070[7:0];
  _RAND_3071 = {1{`RANDOM}};
  lineBuffer_3064 = _RAND_3071[7:0];
  _RAND_3072 = {1{`RANDOM}};
  lineBuffer_3065 = _RAND_3072[7:0];
  _RAND_3073 = {1{`RANDOM}};
  lineBuffer_3066 = _RAND_3073[7:0];
  _RAND_3074 = {1{`RANDOM}};
  lineBuffer_3067 = _RAND_3074[7:0];
  _RAND_3075 = {1{`RANDOM}};
  lineBuffer_3068 = _RAND_3075[7:0];
  _RAND_3076 = {1{`RANDOM}};
  lineBuffer_3069 = _RAND_3076[7:0];
  _RAND_3077 = {1{`RANDOM}};
  lineBuffer_3070 = _RAND_3077[7:0];
  _RAND_3078 = {1{`RANDOM}};
  lineBuffer_3071 = _RAND_3078[7:0];
  _RAND_3079 = {1{`RANDOM}};
  lineBuffer_3072 = _RAND_3079[7:0];
  _RAND_3080 = {1{`RANDOM}};
  lineBuffer_3073 = _RAND_3080[7:0];
  _RAND_3081 = {1{`RANDOM}};
  lineBuffer_3074 = _RAND_3081[7:0];
  _RAND_3082 = {1{`RANDOM}};
  lineBuffer_3075 = _RAND_3082[7:0];
  _RAND_3083 = {1{`RANDOM}};
  lineBuffer_3076 = _RAND_3083[7:0];
  _RAND_3084 = {1{`RANDOM}};
  lineBuffer_3077 = _RAND_3084[7:0];
  _RAND_3085 = {1{`RANDOM}};
  lineBuffer_3078 = _RAND_3085[7:0];
  _RAND_3086 = {1{`RANDOM}};
  lineBuffer_3079 = _RAND_3086[7:0];
  _RAND_3087 = {1{`RANDOM}};
  lineBuffer_3080 = _RAND_3087[7:0];
  _RAND_3088 = {1{`RANDOM}};
  lineBuffer_3081 = _RAND_3088[7:0];
  _RAND_3089 = {1{`RANDOM}};
  lineBuffer_3082 = _RAND_3089[7:0];
  _RAND_3090 = {1{`RANDOM}};
  lineBuffer_3083 = _RAND_3090[7:0];
  _RAND_3091 = {1{`RANDOM}};
  lineBuffer_3084 = _RAND_3091[7:0];
  _RAND_3092 = {1{`RANDOM}};
  lineBuffer_3085 = _RAND_3092[7:0];
  _RAND_3093 = {1{`RANDOM}};
  lineBuffer_3086 = _RAND_3093[7:0];
  _RAND_3094 = {1{`RANDOM}};
  lineBuffer_3087 = _RAND_3094[7:0];
  _RAND_3095 = {1{`RANDOM}};
  lineBuffer_3088 = _RAND_3095[7:0];
  _RAND_3096 = {1{`RANDOM}};
  lineBuffer_3089 = _RAND_3096[7:0];
  _RAND_3097 = {1{`RANDOM}};
  lineBuffer_3090 = _RAND_3097[7:0];
  _RAND_3098 = {1{`RANDOM}};
  lineBuffer_3091 = _RAND_3098[7:0];
  _RAND_3099 = {1{`RANDOM}};
  lineBuffer_3092 = _RAND_3099[7:0];
  _RAND_3100 = {1{`RANDOM}};
  lineBuffer_3093 = _RAND_3100[7:0];
  _RAND_3101 = {1{`RANDOM}};
  lineBuffer_3094 = _RAND_3101[7:0];
  _RAND_3102 = {1{`RANDOM}};
  lineBuffer_3095 = _RAND_3102[7:0];
  _RAND_3103 = {1{`RANDOM}};
  lineBuffer_3096 = _RAND_3103[7:0];
  _RAND_3104 = {1{`RANDOM}};
  lineBuffer_3097 = _RAND_3104[7:0];
  _RAND_3105 = {1{`RANDOM}};
  lineBuffer_3098 = _RAND_3105[7:0];
  _RAND_3106 = {1{`RANDOM}};
  lineBuffer_3099 = _RAND_3106[7:0];
  _RAND_3107 = {1{`RANDOM}};
  lineBuffer_3100 = _RAND_3107[7:0];
  _RAND_3108 = {1{`RANDOM}};
  lineBuffer_3101 = _RAND_3108[7:0];
  _RAND_3109 = {1{`RANDOM}};
  lineBuffer_3102 = _RAND_3109[7:0];
  _RAND_3110 = {1{`RANDOM}};
  lineBuffer_3103 = _RAND_3110[7:0];
  _RAND_3111 = {1{`RANDOM}};
  lineBuffer_3104 = _RAND_3111[7:0];
  _RAND_3112 = {1{`RANDOM}};
  lineBuffer_3105 = _RAND_3112[7:0];
  _RAND_3113 = {1{`RANDOM}};
  lineBuffer_3106 = _RAND_3113[7:0];
  _RAND_3114 = {1{`RANDOM}};
  lineBuffer_3107 = _RAND_3114[7:0];
  _RAND_3115 = {1{`RANDOM}};
  lineBuffer_3108 = _RAND_3115[7:0];
  _RAND_3116 = {1{`RANDOM}};
  lineBuffer_3109 = _RAND_3116[7:0];
  _RAND_3117 = {1{`RANDOM}};
  lineBuffer_3110 = _RAND_3117[7:0];
  _RAND_3118 = {1{`RANDOM}};
  lineBuffer_3111 = _RAND_3118[7:0];
  _RAND_3119 = {1{`RANDOM}};
  lineBuffer_3112 = _RAND_3119[7:0];
  _RAND_3120 = {1{`RANDOM}};
  lineBuffer_3113 = _RAND_3120[7:0];
  _RAND_3121 = {1{`RANDOM}};
  lineBuffer_3114 = _RAND_3121[7:0];
  _RAND_3122 = {1{`RANDOM}};
  lineBuffer_3115 = _RAND_3122[7:0];
  _RAND_3123 = {1{`RANDOM}};
  lineBuffer_3116 = _RAND_3123[7:0];
  _RAND_3124 = {1{`RANDOM}};
  lineBuffer_3117 = _RAND_3124[7:0];
  _RAND_3125 = {1{`RANDOM}};
  lineBuffer_3118 = _RAND_3125[7:0];
  _RAND_3126 = {1{`RANDOM}};
  lineBuffer_3119 = _RAND_3126[7:0];
  _RAND_3127 = {1{`RANDOM}};
  lineBuffer_3120 = _RAND_3127[7:0];
  _RAND_3128 = {1{`RANDOM}};
  lineBuffer_3121 = _RAND_3128[7:0];
  _RAND_3129 = {1{`RANDOM}};
  lineBuffer_3122 = _RAND_3129[7:0];
  _RAND_3130 = {1{`RANDOM}};
  lineBuffer_3123 = _RAND_3130[7:0];
  _RAND_3131 = {1{`RANDOM}};
  lineBuffer_3124 = _RAND_3131[7:0];
  _RAND_3132 = {1{`RANDOM}};
  lineBuffer_3125 = _RAND_3132[7:0];
  _RAND_3133 = {1{`RANDOM}};
  lineBuffer_3126 = _RAND_3133[7:0];
  _RAND_3134 = {1{`RANDOM}};
  lineBuffer_3127 = _RAND_3134[7:0];
  _RAND_3135 = {1{`RANDOM}};
  lineBuffer_3128 = _RAND_3135[7:0];
  _RAND_3136 = {1{`RANDOM}};
  lineBuffer_3129 = _RAND_3136[7:0];
  _RAND_3137 = {1{`RANDOM}};
  lineBuffer_3130 = _RAND_3137[7:0];
  _RAND_3138 = {1{`RANDOM}};
  lineBuffer_3131 = _RAND_3138[7:0];
  _RAND_3139 = {1{`RANDOM}};
  lineBuffer_3132 = _RAND_3139[7:0];
  _RAND_3140 = {1{`RANDOM}};
  lineBuffer_3133 = _RAND_3140[7:0];
  _RAND_3141 = {1{`RANDOM}};
  lineBuffer_3134 = _RAND_3141[7:0];
  _RAND_3142 = {1{`RANDOM}};
  lineBuffer_3135 = _RAND_3142[7:0];
  _RAND_3143 = {1{`RANDOM}};
  lineBuffer_3136 = _RAND_3143[7:0];
  _RAND_3144 = {1{`RANDOM}};
  lineBuffer_3137 = _RAND_3144[7:0];
  _RAND_3145 = {1{`RANDOM}};
  lineBuffer_3138 = _RAND_3145[7:0];
  _RAND_3146 = {1{`RANDOM}};
  lineBuffer_3139 = _RAND_3146[7:0];
  _RAND_3147 = {1{`RANDOM}};
  lineBuffer_3140 = _RAND_3147[7:0];
  _RAND_3148 = {1{`RANDOM}};
  lineBuffer_3141 = _RAND_3148[7:0];
  _RAND_3149 = {1{`RANDOM}};
  lineBuffer_3142 = _RAND_3149[7:0];
  _RAND_3150 = {1{`RANDOM}};
  lineBuffer_3143 = _RAND_3150[7:0];
  _RAND_3151 = {1{`RANDOM}};
  lineBuffer_3144 = _RAND_3151[7:0];
  _RAND_3152 = {1{`RANDOM}};
  lineBuffer_3145 = _RAND_3152[7:0];
  _RAND_3153 = {1{`RANDOM}};
  lineBuffer_3146 = _RAND_3153[7:0];
  _RAND_3154 = {1{`RANDOM}};
  lineBuffer_3147 = _RAND_3154[7:0];
  _RAND_3155 = {1{`RANDOM}};
  lineBuffer_3148 = _RAND_3155[7:0];
  _RAND_3156 = {1{`RANDOM}};
  lineBuffer_3149 = _RAND_3156[7:0];
  _RAND_3157 = {1{`RANDOM}};
  lineBuffer_3150 = _RAND_3157[7:0];
  _RAND_3158 = {1{`RANDOM}};
  lineBuffer_3151 = _RAND_3158[7:0];
  _RAND_3159 = {1{`RANDOM}};
  lineBuffer_3152 = _RAND_3159[7:0];
  _RAND_3160 = {1{`RANDOM}};
  lineBuffer_3153 = _RAND_3160[7:0];
  _RAND_3161 = {1{`RANDOM}};
  lineBuffer_3154 = _RAND_3161[7:0];
  _RAND_3162 = {1{`RANDOM}};
  lineBuffer_3155 = _RAND_3162[7:0];
  _RAND_3163 = {1{`RANDOM}};
  lineBuffer_3156 = _RAND_3163[7:0];
  _RAND_3164 = {1{`RANDOM}};
  lineBuffer_3157 = _RAND_3164[7:0];
  _RAND_3165 = {1{`RANDOM}};
  lineBuffer_3158 = _RAND_3165[7:0];
  _RAND_3166 = {1{`RANDOM}};
  lineBuffer_3159 = _RAND_3166[7:0];
  _RAND_3167 = {1{`RANDOM}};
  lineBuffer_3160 = _RAND_3167[7:0];
  _RAND_3168 = {1{`RANDOM}};
  lineBuffer_3161 = _RAND_3168[7:0];
  _RAND_3169 = {1{`RANDOM}};
  lineBuffer_3162 = _RAND_3169[7:0];
  _RAND_3170 = {1{`RANDOM}};
  lineBuffer_3163 = _RAND_3170[7:0];
  _RAND_3171 = {1{`RANDOM}};
  lineBuffer_3164 = _RAND_3171[7:0];
  _RAND_3172 = {1{`RANDOM}};
  lineBuffer_3165 = _RAND_3172[7:0];
  _RAND_3173 = {1{`RANDOM}};
  lineBuffer_3166 = _RAND_3173[7:0];
  _RAND_3174 = {1{`RANDOM}};
  lineBuffer_3167 = _RAND_3174[7:0];
  _RAND_3175 = {1{`RANDOM}};
  lineBuffer_3168 = _RAND_3175[7:0];
  _RAND_3176 = {1{`RANDOM}};
  lineBuffer_3169 = _RAND_3176[7:0];
  _RAND_3177 = {1{`RANDOM}};
  lineBuffer_3170 = _RAND_3177[7:0];
  _RAND_3178 = {1{`RANDOM}};
  lineBuffer_3171 = _RAND_3178[7:0];
  _RAND_3179 = {1{`RANDOM}};
  lineBuffer_3172 = _RAND_3179[7:0];
  _RAND_3180 = {1{`RANDOM}};
  lineBuffer_3173 = _RAND_3180[7:0];
  _RAND_3181 = {1{`RANDOM}};
  lineBuffer_3174 = _RAND_3181[7:0];
  _RAND_3182 = {1{`RANDOM}};
  lineBuffer_3175 = _RAND_3182[7:0];
  _RAND_3183 = {1{`RANDOM}};
  lineBuffer_3176 = _RAND_3183[7:0];
  _RAND_3184 = {1{`RANDOM}};
  lineBuffer_3177 = _RAND_3184[7:0];
  _RAND_3185 = {1{`RANDOM}};
  lineBuffer_3178 = _RAND_3185[7:0];
  _RAND_3186 = {1{`RANDOM}};
  lineBuffer_3179 = _RAND_3186[7:0];
  _RAND_3187 = {1{`RANDOM}};
  lineBuffer_3180 = _RAND_3187[7:0];
  _RAND_3188 = {1{`RANDOM}};
  lineBuffer_3181 = _RAND_3188[7:0];
  _RAND_3189 = {1{`RANDOM}};
  lineBuffer_3182 = _RAND_3189[7:0];
  _RAND_3190 = {1{`RANDOM}};
  lineBuffer_3183 = _RAND_3190[7:0];
  _RAND_3191 = {1{`RANDOM}};
  lineBuffer_3184 = _RAND_3191[7:0];
  _RAND_3192 = {1{`RANDOM}};
  lineBuffer_3185 = _RAND_3192[7:0];
  _RAND_3193 = {1{`RANDOM}};
  lineBuffer_3186 = _RAND_3193[7:0];
  _RAND_3194 = {1{`RANDOM}};
  lineBuffer_3187 = _RAND_3194[7:0];
  _RAND_3195 = {1{`RANDOM}};
  lineBuffer_3188 = _RAND_3195[7:0];
  _RAND_3196 = {1{`RANDOM}};
  lineBuffer_3189 = _RAND_3196[7:0];
  _RAND_3197 = {1{`RANDOM}};
  lineBuffer_3190 = _RAND_3197[7:0];
  _RAND_3198 = {1{`RANDOM}};
  lineBuffer_3191 = _RAND_3198[7:0];
  _RAND_3199 = {1{`RANDOM}};
  lineBuffer_3192 = _RAND_3199[7:0];
  _RAND_3200 = {1{`RANDOM}};
  lineBuffer_3193 = _RAND_3200[7:0];
  _RAND_3201 = {1{`RANDOM}};
  lineBuffer_3194 = _RAND_3201[7:0];
  _RAND_3202 = {1{`RANDOM}};
  lineBuffer_3195 = _RAND_3202[7:0];
  _RAND_3203 = {1{`RANDOM}};
  lineBuffer_3196 = _RAND_3203[7:0];
  _RAND_3204 = {1{`RANDOM}};
  lineBuffer_3197 = _RAND_3204[7:0];
  _RAND_3205 = {1{`RANDOM}};
  lineBuffer_3198 = _RAND_3205[7:0];
  _RAND_3206 = {1{`RANDOM}};
  lineBuffer_3199 = _RAND_3206[7:0];
  _RAND_3207 = {1{`RANDOM}};
  lineBuffer_3200 = _RAND_3207[7:0];
  _RAND_3208 = {1{`RANDOM}};
  lineBuffer_3201 = _RAND_3208[7:0];
  _RAND_3209 = {1{`RANDOM}};
  lineBuffer_3202 = _RAND_3209[7:0];
  _RAND_3210 = {1{`RANDOM}};
  lineBuffer_3203 = _RAND_3210[7:0];
  _RAND_3211 = {1{`RANDOM}};
  lineBuffer_3204 = _RAND_3211[7:0];
  _RAND_3212 = {1{`RANDOM}};
  lineBuffer_3205 = _RAND_3212[7:0];
  _RAND_3213 = {1{`RANDOM}};
  lineBuffer_3206 = _RAND_3213[7:0];
  _RAND_3214 = {1{`RANDOM}};
  lineBuffer_3207 = _RAND_3214[7:0];
  _RAND_3215 = {1{`RANDOM}};
  lineBuffer_3208 = _RAND_3215[7:0];
  _RAND_3216 = {1{`RANDOM}};
  lineBuffer_3209 = _RAND_3216[7:0];
  _RAND_3217 = {1{`RANDOM}};
  lineBuffer_3210 = _RAND_3217[7:0];
  _RAND_3218 = {1{`RANDOM}};
  lineBuffer_3211 = _RAND_3218[7:0];
  _RAND_3219 = {1{`RANDOM}};
  lineBuffer_3212 = _RAND_3219[7:0];
  _RAND_3220 = {1{`RANDOM}};
  lineBuffer_3213 = _RAND_3220[7:0];
  _RAND_3221 = {1{`RANDOM}};
  lineBuffer_3214 = _RAND_3221[7:0];
  _RAND_3222 = {1{`RANDOM}};
  lineBuffer_3215 = _RAND_3222[7:0];
  _RAND_3223 = {1{`RANDOM}};
  lineBuffer_3216 = _RAND_3223[7:0];
  _RAND_3224 = {1{`RANDOM}};
  lineBuffer_3217 = _RAND_3224[7:0];
  _RAND_3225 = {1{`RANDOM}};
  lineBuffer_3218 = _RAND_3225[7:0];
  _RAND_3226 = {1{`RANDOM}};
  lineBuffer_3219 = _RAND_3226[7:0];
  _RAND_3227 = {1{`RANDOM}};
  lineBuffer_3220 = _RAND_3227[7:0];
  _RAND_3228 = {1{`RANDOM}};
  lineBuffer_3221 = _RAND_3228[7:0];
  _RAND_3229 = {1{`RANDOM}};
  lineBuffer_3222 = _RAND_3229[7:0];
  _RAND_3230 = {1{`RANDOM}};
  lineBuffer_3223 = _RAND_3230[7:0];
  _RAND_3231 = {1{`RANDOM}};
  lineBuffer_3224 = _RAND_3231[7:0];
  _RAND_3232 = {1{`RANDOM}};
  lineBuffer_3225 = _RAND_3232[7:0];
  _RAND_3233 = {1{`RANDOM}};
  lineBuffer_3226 = _RAND_3233[7:0];
  _RAND_3234 = {1{`RANDOM}};
  lineBuffer_3227 = _RAND_3234[7:0];
  _RAND_3235 = {1{`RANDOM}};
  lineBuffer_3228 = _RAND_3235[7:0];
  _RAND_3236 = {1{`RANDOM}};
  lineBuffer_3229 = _RAND_3236[7:0];
  _RAND_3237 = {1{`RANDOM}};
  lineBuffer_3230 = _RAND_3237[7:0];
  _RAND_3238 = {1{`RANDOM}};
  lineBuffer_3231 = _RAND_3238[7:0];
  _RAND_3239 = {1{`RANDOM}};
  lineBuffer_3232 = _RAND_3239[7:0];
  _RAND_3240 = {1{`RANDOM}};
  lineBuffer_3233 = _RAND_3240[7:0];
  _RAND_3241 = {1{`RANDOM}};
  lineBuffer_3234 = _RAND_3241[7:0];
  _RAND_3242 = {1{`RANDOM}};
  lineBuffer_3235 = _RAND_3242[7:0];
  _RAND_3243 = {1{`RANDOM}};
  lineBuffer_3236 = _RAND_3243[7:0];
  _RAND_3244 = {1{`RANDOM}};
  lineBuffer_3237 = _RAND_3244[7:0];
  _RAND_3245 = {1{`RANDOM}};
  lineBuffer_3238 = _RAND_3245[7:0];
  _RAND_3246 = {1{`RANDOM}};
  lineBuffer_3239 = _RAND_3246[7:0];
  _RAND_3247 = {1{`RANDOM}};
  lineBuffer_3240 = _RAND_3247[7:0];
  _RAND_3248 = {1{`RANDOM}};
  lineBuffer_3241 = _RAND_3248[7:0];
  _RAND_3249 = {1{`RANDOM}};
  lineBuffer_3242 = _RAND_3249[7:0];
  _RAND_3250 = {1{`RANDOM}};
  lineBuffer_3243 = _RAND_3250[7:0];
  _RAND_3251 = {1{`RANDOM}};
  lineBuffer_3244 = _RAND_3251[7:0];
  _RAND_3252 = {1{`RANDOM}};
  lineBuffer_3245 = _RAND_3252[7:0];
  _RAND_3253 = {1{`RANDOM}};
  lineBuffer_3246 = _RAND_3253[7:0];
  _RAND_3254 = {1{`RANDOM}};
  lineBuffer_3247 = _RAND_3254[7:0];
  _RAND_3255 = {1{`RANDOM}};
  lineBuffer_3248 = _RAND_3255[7:0];
  _RAND_3256 = {1{`RANDOM}};
  lineBuffer_3249 = _RAND_3256[7:0];
  _RAND_3257 = {1{`RANDOM}};
  lineBuffer_3250 = _RAND_3257[7:0];
  _RAND_3258 = {1{`RANDOM}};
  lineBuffer_3251 = _RAND_3258[7:0];
  _RAND_3259 = {1{`RANDOM}};
  lineBuffer_3252 = _RAND_3259[7:0];
  _RAND_3260 = {1{`RANDOM}};
  lineBuffer_3253 = _RAND_3260[7:0];
  _RAND_3261 = {1{`RANDOM}};
  lineBuffer_3254 = _RAND_3261[7:0];
  _RAND_3262 = {1{`RANDOM}};
  lineBuffer_3255 = _RAND_3262[7:0];
  _RAND_3263 = {1{`RANDOM}};
  lineBuffer_3256 = _RAND_3263[7:0];
  _RAND_3264 = {1{`RANDOM}};
  lineBuffer_3257 = _RAND_3264[7:0];
  _RAND_3265 = {1{`RANDOM}};
  lineBuffer_3258 = _RAND_3265[7:0];
  _RAND_3266 = {1{`RANDOM}};
  lineBuffer_3259 = _RAND_3266[7:0];
  _RAND_3267 = {1{`RANDOM}};
  lineBuffer_3260 = _RAND_3267[7:0];
  _RAND_3268 = {1{`RANDOM}};
  lineBuffer_3261 = _RAND_3268[7:0];
  _RAND_3269 = {1{`RANDOM}};
  lineBuffer_3262 = _RAND_3269[7:0];
  _RAND_3270 = {1{`RANDOM}};
  lineBuffer_3263 = _RAND_3270[7:0];
  _RAND_3271 = {1{`RANDOM}};
  lineBuffer_3264 = _RAND_3271[7:0];
  _RAND_3272 = {1{`RANDOM}};
  lineBuffer_3265 = _RAND_3272[7:0];
  _RAND_3273 = {1{`RANDOM}};
  lineBuffer_3266 = _RAND_3273[7:0];
  _RAND_3274 = {1{`RANDOM}};
  lineBuffer_3267 = _RAND_3274[7:0];
  _RAND_3275 = {1{`RANDOM}};
  lineBuffer_3268 = _RAND_3275[7:0];
  _RAND_3276 = {1{`RANDOM}};
  lineBuffer_3269 = _RAND_3276[7:0];
  _RAND_3277 = {1{`RANDOM}};
  lineBuffer_3270 = _RAND_3277[7:0];
  _RAND_3278 = {1{`RANDOM}};
  lineBuffer_3271 = _RAND_3278[7:0];
  _RAND_3279 = {1{`RANDOM}};
  lineBuffer_3272 = _RAND_3279[7:0];
  _RAND_3280 = {1{`RANDOM}};
  lineBuffer_3273 = _RAND_3280[7:0];
  _RAND_3281 = {1{`RANDOM}};
  lineBuffer_3274 = _RAND_3281[7:0];
  _RAND_3282 = {1{`RANDOM}};
  lineBuffer_3275 = _RAND_3282[7:0];
  _RAND_3283 = {1{`RANDOM}};
  lineBuffer_3276 = _RAND_3283[7:0];
  _RAND_3284 = {1{`RANDOM}};
  lineBuffer_3277 = _RAND_3284[7:0];
  _RAND_3285 = {1{`RANDOM}};
  lineBuffer_3278 = _RAND_3285[7:0];
  _RAND_3286 = {1{`RANDOM}};
  lineBuffer_3279 = _RAND_3286[7:0];
  _RAND_3287 = {1{`RANDOM}};
  lineBuffer_3280 = _RAND_3287[7:0];
  _RAND_3288 = {1{`RANDOM}};
  lineBuffer_3281 = _RAND_3288[7:0];
  _RAND_3289 = {1{`RANDOM}};
  lineBuffer_3282 = _RAND_3289[7:0];
  _RAND_3290 = {1{`RANDOM}};
  lineBuffer_3283 = _RAND_3290[7:0];
  _RAND_3291 = {1{`RANDOM}};
  lineBuffer_3284 = _RAND_3291[7:0];
  _RAND_3292 = {1{`RANDOM}};
  lineBuffer_3285 = _RAND_3292[7:0];
  _RAND_3293 = {1{`RANDOM}};
  lineBuffer_3286 = _RAND_3293[7:0];
  _RAND_3294 = {1{`RANDOM}};
  lineBuffer_3287 = _RAND_3294[7:0];
  _RAND_3295 = {1{`RANDOM}};
  lineBuffer_3288 = _RAND_3295[7:0];
  _RAND_3296 = {1{`RANDOM}};
  lineBuffer_3289 = _RAND_3296[7:0];
  _RAND_3297 = {1{`RANDOM}};
  lineBuffer_3290 = _RAND_3297[7:0];
  _RAND_3298 = {1{`RANDOM}};
  lineBuffer_3291 = _RAND_3298[7:0];
  _RAND_3299 = {1{`RANDOM}};
  lineBuffer_3292 = _RAND_3299[7:0];
  _RAND_3300 = {1{`RANDOM}};
  lineBuffer_3293 = _RAND_3300[7:0];
  _RAND_3301 = {1{`RANDOM}};
  lineBuffer_3294 = _RAND_3301[7:0];
  _RAND_3302 = {1{`RANDOM}};
  lineBuffer_3295 = _RAND_3302[7:0];
  _RAND_3303 = {1{`RANDOM}};
  lineBuffer_3296 = _RAND_3303[7:0];
  _RAND_3304 = {1{`RANDOM}};
  lineBuffer_3297 = _RAND_3304[7:0];
  _RAND_3305 = {1{`RANDOM}};
  lineBuffer_3298 = _RAND_3305[7:0];
  _RAND_3306 = {1{`RANDOM}};
  lineBuffer_3299 = _RAND_3306[7:0];
  _RAND_3307 = {1{`RANDOM}};
  lineBuffer_3300 = _RAND_3307[7:0];
  _RAND_3308 = {1{`RANDOM}};
  lineBuffer_3301 = _RAND_3308[7:0];
  _RAND_3309 = {1{`RANDOM}};
  lineBuffer_3302 = _RAND_3309[7:0];
  _RAND_3310 = {1{`RANDOM}};
  lineBuffer_3303 = _RAND_3310[7:0];
  _RAND_3311 = {1{`RANDOM}};
  lineBuffer_3304 = _RAND_3311[7:0];
  _RAND_3312 = {1{`RANDOM}};
  lineBuffer_3305 = _RAND_3312[7:0];
  _RAND_3313 = {1{`RANDOM}};
  lineBuffer_3306 = _RAND_3313[7:0];
  _RAND_3314 = {1{`RANDOM}};
  lineBuffer_3307 = _RAND_3314[7:0];
  _RAND_3315 = {1{`RANDOM}};
  lineBuffer_3308 = _RAND_3315[7:0];
  _RAND_3316 = {1{`RANDOM}};
  lineBuffer_3309 = _RAND_3316[7:0];
  _RAND_3317 = {1{`RANDOM}};
  lineBuffer_3310 = _RAND_3317[7:0];
  _RAND_3318 = {1{`RANDOM}};
  lineBuffer_3311 = _RAND_3318[7:0];
  _RAND_3319 = {1{`RANDOM}};
  lineBuffer_3312 = _RAND_3319[7:0];
  _RAND_3320 = {1{`RANDOM}};
  lineBuffer_3313 = _RAND_3320[7:0];
  _RAND_3321 = {1{`RANDOM}};
  lineBuffer_3314 = _RAND_3321[7:0];
  _RAND_3322 = {1{`RANDOM}};
  lineBuffer_3315 = _RAND_3322[7:0];
  _RAND_3323 = {1{`RANDOM}};
  lineBuffer_3316 = _RAND_3323[7:0];
  _RAND_3324 = {1{`RANDOM}};
  lineBuffer_3317 = _RAND_3324[7:0];
  _RAND_3325 = {1{`RANDOM}};
  lineBuffer_3318 = _RAND_3325[7:0];
  _RAND_3326 = {1{`RANDOM}};
  lineBuffer_3319 = _RAND_3326[7:0];
  _RAND_3327 = {1{`RANDOM}};
  lineBuffer_3320 = _RAND_3327[7:0];
  _RAND_3328 = {1{`RANDOM}};
  lineBuffer_3321 = _RAND_3328[7:0];
  _RAND_3329 = {1{`RANDOM}};
  lineBuffer_3322 = _RAND_3329[7:0];
  _RAND_3330 = {1{`RANDOM}};
  lineBuffer_3323 = _RAND_3330[7:0];
  _RAND_3331 = {1{`RANDOM}};
  lineBuffer_3324 = _RAND_3331[7:0];
  _RAND_3332 = {1{`RANDOM}};
  lineBuffer_3325 = _RAND_3332[7:0];
  _RAND_3333 = {1{`RANDOM}};
  lineBuffer_3326 = _RAND_3333[7:0];
  _RAND_3334 = {1{`RANDOM}};
  lineBuffer_3327 = _RAND_3334[7:0];
  _RAND_3335 = {1{`RANDOM}};
  lineBuffer_3328 = _RAND_3335[7:0];
  _RAND_3336 = {1{`RANDOM}};
  lineBuffer_3329 = _RAND_3336[7:0];
  _RAND_3337 = {1{`RANDOM}};
  lineBuffer_3330 = _RAND_3337[7:0];
  _RAND_3338 = {1{`RANDOM}};
  lineBuffer_3331 = _RAND_3338[7:0];
  _RAND_3339 = {1{`RANDOM}};
  lineBuffer_3332 = _RAND_3339[7:0];
  _RAND_3340 = {1{`RANDOM}};
  lineBuffer_3333 = _RAND_3340[7:0];
  _RAND_3341 = {1{`RANDOM}};
  lineBuffer_3334 = _RAND_3341[7:0];
  _RAND_3342 = {1{`RANDOM}};
  lineBuffer_3335 = _RAND_3342[7:0];
  _RAND_3343 = {1{`RANDOM}};
  lineBuffer_3336 = _RAND_3343[7:0];
  _RAND_3344 = {1{`RANDOM}};
  lineBuffer_3337 = _RAND_3344[7:0];
  _RAND_3345 = {1{`RANDOM}};
  lineBuffer_3338 = _RAND_3345[7:0];
  _RAND_3346 = {1{`RANDOM}};
  lineBuffer_3339 = _RAND_3346[7:0];
  _RAND_3347 = {1{`RANDOM}};
  lineBuffer_3340 = _RAND_3347[7:0];
  _RAND_3348 = {1{`RANDOM}};
  lineBuffer_3341 = _RAND_3348[7:0];
  _RAND_3349 = {1{`RANDOM}};
  lineBuffer_3342 = _RAND_3349[7:0];
  _RAND_3350 = {1{`RANDOM}};
  lineBuffer_3343 = _RAND_3350[7:0];
  _RAND_3351 = {1{`RANDOM}};
  lineBuffer_3344 = _RAND_3351[7:0];
  _RAND_3352 = {1{`RANDOM}};
  lineBuffer_3345 = _RAND_3352[7:0];
  _RAND_3353 = {1{`RANDOM}};
  lineBuffer_3346 = _RAND_3353[7:0];
  _RAND_3354 = {1{`RANDOM}};
  lineBuffer_3347 = _RAND_3354[7:0];
  _RAND_3355 = {1{`RANDOM}};
  lineBuffer_3348 = _RAND_3355[7:0];
  _RAND_3356 = {1{`RANDOM}};
  lineBuffer_3349 = _RAND_3356[7:0];
  _RAND_3357 = {1{`RANDOM}};
  lineBuffer_3350 = _RAND_3357[7:0];
  _RAND_3358 = {1{`RANDOM}};
  lineBuffer_3351 = _RAND_3358[7:0];
  _RAND_3359 = {1{`RANDOM}};
  lineBuffer_3352 = _RAND_3359[7:0];
  _RAND_3360 = {1{`RANDOM}};
  lineBuffer_3353 = _RAND_3360[7:0];
  _RAND_3361 = {1{`RANDOM}};
  lineBuffer_3354 = _RAND_3361[7:0];
  _RAND_3362 = {1{`RANDOM}};
  lineBuffer_3355 = _RAND_3362[7:0];
  _RAND_3363 = {1{`RANDOM}};
  lineBuffer_3356 = _RAND_3363[7:0];
  _RAND_3364 = {1{`RANDOM}};
  lineBuffer_3357 = _RAND_3364[7:0];
  _RAND_3365 = {1{`RANDOM}};
  lineBuffer_3358 = _RAND_3365[7:0];
  _RAND_3366 = {1{`RANDOM}};
  lineBuffer_3359 = _RAND_3366[7:0];
  _RAND_3367 = {1{`RANDOM}};
  lineBuffer_3360 = _RAND_3367[7:0];
  _RAND_3368 = {1{`RANDOM}};
  lineBuffer_3361 = _RAND_3368[7:0];
  _RAND_3369 = {1{`RANDOM}};
  lineBuffer_3362 = _RAND_3369[7:0];
  _RAND_3370 = {1{`RANDOM}};
  lineBuffer_3363 = _RAND_3370[7:0];
  _RAND_3371 = {1{`RANDOM}};
  lineBuffer_3364 = _RAND_3371[7:0];
  _RAND_3372 = {1{`RANDOM}};
  lineBuffer_3365 = _RAND_3372[7:0];
  _RAND_3373 = {1{`RANDOM}};
  lineBuffer_3366 = _RAND_3373[7:0];
  _RAND_3374 = {1{`RANDOM}};
  lineBuffer_3367 = _RAND_3374[7:0];
  _RAND_3375 = {1{`RANDOM}};
  lineBuffer_3368 = _RAND_3375[7:0];
  _RAND_3376 = {1{`RANDOM}};
  lineBuffer_3369 = _RAND_3376[7:0];
  _RAND_3377 = {1{`RANDOM}};
  lineBuffer_3370 = _RAND_3377[7:0];
  _RAND_3378 = {1{`RANDOM}};
  lineBuffer_3371 = _RAND_3378[7:0];
  _RAND_3379 = {1{`RANDOM}};
  lineBuffer_3372 = _RAND_3379[7:0];
  _RAND_3380 = {1{`RANDOM}};
  lineBuffer_3373 = _RAND_3380[7:0];
  _RAND_3381 = {1{`RANDOM}};
  lineBuffer_3374 = _RAND_3381[7:0];
  _RAND_3382 = {1{`RANDOM}};
  lineBuffer_3375 = _RAND_3382[7:0];
  _RAND_3383 = {1{`RANDOM}};
  lineBuffer_3376 = _RAND_3383[7:0];
  _RAND_3384 = {1{`RANDOM}};
  lineBuffer_3377 = _RAND_3384[7:0];
  _RAND_3385 = {1{`RANDOM}};
  lineBuffer_3378 = _RAND_3385[7:0];
  _RAND_3386 = {1{`RANDOM}};
  lineBuffer_3379 = _RAND_3386[7:0];
  _RAND_3387 = {1{`RANDOM}};
  lineBuffer_3380 = _RAND_3387[7:0];
  _RAND_3388 = {1{`RANDOM}};
  lineBuffer_3381 = _RAND_3388[7:0];
  _RAND_3389 = {1{`RANDOM}};
  lineBuffer_3382 = _RAND_3389[7:0];
  _RAND_3390 = {1{`RANDOM}};
  lineBuffer_3383 = _RAND_3390[7:0];
  _RAND_3391 = {1{`RANDOM}};
  lineBuffer_3384 = _RAND_3391[7:0];
  _RAND_3392 = {1{`RANDOM}};
  lineBuffer_3385 = _RAND_3392[7:0];
  _RAND_3393 = {1{`RANDOM}};
  lineBuffer_3386 = _RAND_3393[7:0];
  _RAND_3394 = {1{`RANDOM}};
  lineBuffer_3387 = _RAND_3394[7:0];
  _RAND_3395 = {1{`RANDOM}};
  lineBuffer_3388 = _RAND_3395[7:0];
  _RAND_3396 = {1{`RANDOM}};
  lineBuffer_3389 = _RAND_3396[7:0];
  _RAND_3397 = {1{`RANDOM}};
  lineBuffer_3390 = _RAND_3397[7:0];
  _RAND_3398 = {1{`RANDOM}};
  lineBuffer_3391 = _RAND_3398[7:0];
  _RAND_3399 = {1{`RANDOM}};
  lineBuffer_3392 = _RAND_3399[7:0];
  _RAND_3400 = {1{`RANDOM}};
  lineBuffer_3393 = _RAND_3400[7:0];
  _RAND_3401 = {1{`RANDOM}};
  lineBuffer_3394 = _RAND_3401[7:0];
  _RAND_3402 = {1{`RANDOM}};
  lineBuffer_3395 = _RAND_3402[7:0];
  _RAND_3403 = {1{`RANDOM}};
  lineBuffer_3396 = _RAND_3403[7:0];
  _RAND_3404 = {1{`RANDOM}};
  lineBuffer_3397 = _RAND_3404[7:0];
  _RAND_3405 = {1{`RANDOM}};
  lineBuffer_3398 = _RAND_3405[7:0];
  _RAND_3406 = {1{`RANDOM}};
  lineBuffer_3399 = _RAND_3406[7:0];
  _RAND_3407 = {1{`RANDOM}};
  lineBuffer_3400 = _RAND_3407[7:0];
  _RAND_3408 = {1{`RANDOM}};
  lineBuffer_3401 = _RAND_3408[7:0];
  _RAND_3409 = {1{`RANDOM}};
  lineBuffer_3402 = _RAND_3409[7:0];
  _RAND_3410 = {1{`RANDOM}};
  lineBuffer_3403 = _RAND_3410[7:0];
  _RAND_3411 = {1{`RANDOM}};
  lineBuffer_3404 = _RAND_3411[7:0];
  _RAND_3412 = {1{`RANDOM}};
  lineBuffer_3405 = _RAND_3412[7:0];
  _RAND_3413 = {1{`RANDOM}};
  lineBuffer_3406 = _RAND_3413[7:0];
  _RAND_3414 = {1{`RANDOM}};
  lineBuffer_3407 = _RAND_3414[7:0];
  _RAND_3415 = {1{`RANDOM}};
  lineBuffer_3408 = _RAND_3415[7:0];
  _RAND_3416 = {1{`RANDOM}};
  lineBuffer_3409 = _RAND_3416[7:0];
  _RAND_3417 = {1{`RANDOM}};
  lineBuffer_3410 = _RAND_3417[7:0];
  _RAND_3418 = {1{`RANDOM}};
  lineBuffer_3411 = _RAND_3418[7:0];
  _RAND_3419 = {1{`RANDOM}};
  lineBuffer_3412 = _RAND_3419[7:0];
  _RAND_3420 = {1{`RANDOM}};
  lineBuffer_3413 = _RAND_3420[7:0];
  _RAND_3421 = {1{`RANDOM}};
  lineBuffer_3414 = _RAND_3421[7:0];
  _RAND_3422 = {1{`RANDOM}};
  lineBuffer_3415 = _RAND_3422[7:0];
  _RAND_3423 = {1{`RANDOM}};
  lineBuffer_3416 = _RAND_3423[7:0];
  _RAND_3424 = {1{`RANDOM}};
  lineBuffer_3417 = _RAND_3424[7:0];
  _RAND_3425 = {1{`RANDOM}};
  lineBuffer_3418 = _RAND_3425[7:0];
  _RAND_3426 = {1{`RANDOM}};
  lineBuffer_3419 = _RAND_3426[7:0];
  _RAND_3427 = {1{`RANDOM}};
  lineBuffer_3420 = _RAND_3427[7:0];
  _RAND_3428 = {1{`RANDOM}};
  lineBuffer_3421 = _RAND_3428[7:0];
  _RAND_3429 = {1{`RANDOM}};
  lineBuffer_3422 = _RAND_3429[7:0];
  _RAND_3430 = {1{`RANDOM}};
  lineBuffer_3423 = _RAND_3430[7:0];
  _RAND_3431 = {1{`RANDOM}};
  lineBuffer_3424 = _RAND_3431[7:0];
  _RAND_3432 = {1{`RANDOM}};
  lineBuffer_3425 = _RAND_3432[7:0];
  _RAND_3433 = {1{`RANDOM}};
  lineBuffer_3426 = _RAND_3433[7:0];
  _RAND_3434 = {1{`RANDOM}};
  lineBuffer_3427 = _RAND_3434[7:0];
  _RAND_3435 = {1{`RANDOM}};
  lineBuffer_3428 = _RAND_3435[7:0];
  _RAND_3436 = {1{`RANDOM}};
  lineBuffer_3429 = _RAND_3436[7:0];
  _RAND_3437 = {1{`RANDOM}};
  lineBuffer_3430 = _RAND_3437[7:0];
  _RAND_3438 = {1{`RANDOM}};
  lineBuffer_3431 = _RAND_3438[7:0];
  _RAND_3439 = {1{`RANDOM}};
  lineBuffer_3432 = _RAND_3439[7:0];
  _RAND_3440 = {1{`RANDOM}};
  lineBuffer_3433 = _RAND_3440[7:0];
  _RAND_3441 = {1{`RANDOM}};
  lineBuffer_3434 = _RAND_3441[7:0];
  _RAND_3442 = {1{`RANDOM}};
  lineBuffer_3435 = _RAND_3442[7:0];
  _RAND_3443 = {1{`RANDOM}};
  lineBuffer_3436 = _RAND_3443[7:0];
  _RAND_3444 = {1{`RANDOM}};
  lineBuffer_3437 = _RAND_3444[7:0];
  _RAND_3445 = {1{`RANDOM}};
  lineBuffer_3438 = _RAND_3445[7:0];
  _RAND_3446 = {1{`RANDOM}};
  lineBuffer_3439 = _RAND_3446[7:0];
  _RAND_3447 = {1{`RANDOM}};
  lineBuffer_3440 = _RAND_3447[7:0];
  _RAND_3448 = {1{`RANDOM}};
  lineBuffer_3441 = _RAND_3448[7:0];
  _RAND_3449 = {1{`RANDOM}};
  lineBuffer_3442 = _RAND_3449[7:0];
  _RAND_3450 = {1{`RANDOM}};
  lineBuffer_3443 = _RAND_3450[7:0];
  _RAND_3451 = {1{`RANDOM}};
  lineBuffer_3444 = _RAND_3451[7:0];
  _RAND_3452 = {1{`RANDOM}};
  lineBuffer_3445 = _RAND_3452[7:0];
  _RAND_3453 = {1{`RANDOM}};
  lineBuffer_3446 = _RAND_3453[7:0];
  _RAND_3454 = {1{`RANDOM}};
  lineBuffer_3447 = _RAND_3454[7:0];
  _RAND_3455 = {1{`RANDOM}};
  lineBuffer_3448 = _RAND_3455[7:0];
  _RAND_3456 = {1{`RANDOM}};
  lineBuffer_3449 = _RAND_3456[7:0];
  _RAND_3457 = {1{`RANDOM}};
  lineBuffer_3450 = _RAND_3457[7:0];
  _RAND_3458 = {1{`RANDOM}};
  lineBuffer_3451 = _RAND_3458[7:0];
  _RAND_3459 = {1{`RANDOM}};
  lineBuffer_3452 = _RAND_3459[7:0];
  _RAND_3460 = {1{`RANDOM}};
  lineBuffer_3453 = _RAND_3460[7:0];
  _RAND_3461 = {1{`RANDOM}};
  lineBuffer_3454 = _RAND_3461[7:0];
  _RAND_3462 = {1{`RANDOM}};
  lineBuffer_3455 = _RAND_3462[7:0];
  _RAND_3463 = {1{`RANDOM}};
  lineBuffer_3456 = _RAND_3463[7:0];
  _RAND_3464 = {1{`RANDOM}};
  lineBuffer_3457 = _RAND_3464[7:0];
  _RAND_3465 = {1{`RANDOM}};
  lineBuffer_3458 = _RAND_3465[7:0];
  _RAND_3466 = {1{`RANDOM}};
  lineBuffer_3459 = _RAND_3466[7:0];
  _RAND_3467 = {1{`RANDOM}};
  lineBuffer_3460 = _RAND_3467[7:0];
  _RAND_3468 = {1{`RANDOM}};
  lineBuffer_3461 = _RAND_3468[7:0];
  _RAND_3469 = {1{`RANDOM}};
  lineBuffer_3462 = _RAND_3469[7:0];
  _RAND_3470 = {1{`RANDOM}};
  lineBuffer_3463 = _RAND_3470[7:0];
  _RAND_3471 = {1{`RANDOM}};
  lineBuffer_3464 = _RAND_3471[7:0];
  _RAND_3472 = {1{`RANDOM}};
  lineBuffer_3465 = _RAND_3472[7:0];
  _RAND_3473 = {1{`RANDOM}};
  lineBuffer_3466 = _RAND_3473[7:0];
  _RAND_3474 = {1{`RANDOM}};
  lineBuffer_3467 = _RAND_3474[7:0];
  _RAND_3475 = {1{`RANDOM}};
  lineBuffer_3468 = _RAND_3475[7:0];
  _RAND_3476 = {1{`RANDOM}};
  lineBuffer_3469 = _RAND_3476[7:0];
  _RAND_3477 = {1{`RANDOM}};
  lineBuffer_3470 = _RAND_3477[7:0];
  _RAND_3478 = {1{`RANDOM}};
  lineBuffer_3471 = _RAND_3478[7:0];
  _RAND_3479 = {1{`RANDOM}};
  lineBuffer_3472 = _RAND_3479[7:0];
  _RAND_3480 = {1{`RANDOM}};
  lineBuffer_3473 = _RAND_3480[7:0];
  _RAND_3481 = {1{`RANDOM}};
  lineBuffer_3474 = _RAND_3481[7:0];
  _RAND_3482 = {1{`RANDOM}};
  lineBuffer_3475 = _RAND_3482[7:0];
  _RAND_3483 = {1{`RANDOM}};
  lineBuffer_3476 = _RAND_3483[7:0];
  _RAND_3484 = {1{`RANDOM}};
  lineBuffer_3477 = _RAND_3484[7:0];
  _RAND_3485 = {1{`RANDOM}};
  lineBuffer_3478 = _RAND_3485[7:0];
  _RAND_3486 = {1{`RANDOM}};
  lineBuffer_3479 = _RAND_3486[7:0];
  _RAND_3487 = {1{`RANDOM}};
  lineBuffer_3480 = _RAND_3487[7:0];
  _RAND_3488 = {1{`RANDOM}};
  lineBuffer_3481 = _RAND_3488[7:0];
  _RAND_3489 = {1{`RANDOM}};
  lineBuffer_3482 = _RAND_3489[7:0];
  _RAND_3490 = {1{`RANDOM}};
  lineBuffer_3483 = _RAND_3490[7:0];
  _RAND_3491 = {1{`RANDOM}};
  lineBuffer_3484 = _RAND_3491[7:0];
  _RAND_3492 = {1{`RANDOM}};
  lineBuffer_3485 = _RAND_3492[7:0];
  _RAND_3493 = {1{`RANDOM}};
  lineBuffer_3486 = _RAND_3493[7:0];
  _RAND_3494 = {1{`RANDOM}};
  lineBuffer_3487 = _RAND_3494[7:0];
  _RAND_3495 = {1{`RANDOM}};
  lineBuffer_3488 = _RAND_3495[7:0];
  _RAND_3496 = {1{`RANDOM}};
  lineBuffer_3489 = _RAND_3496[7:0];
  _RAND_3497 = {1{`RANDOM}};
  lineBuffer_3490 = _RAND_3497[7:0];
  _RAND_3498 = {1{`RANDOM}};
  lineBuffer_3491 = _RAND_3498[7:0];
  _RAND_3499 = {1{`RANDOM}};
  lineBuffer_3492 = _RAND_3499[7:0];
  _RAND_3500 = {1{`RANDOM}};
  lineBuffer_3493 = _RAND_3500[7:0];
  _RAND_3501 = {1{`RANDOM}};
  lineBuffer_3494 = _RAND_3501[7:0];
  _RAND_3502 = {1{`RANDOM}};
  lineBuffer_3495 = _RAND_3502[7:0];
  _RAND_3503 = {1{`RANDOM}};
  lineBuffer_3496 = _RAND_3503[7:0];
  _RAND_3504 = {1{`RANDOM}};
  lineBuffer_3497 = _RAND_3504[7:0];
  _RAND_3505 = {1{`RANDOM}};
  lineBuffer_3498 = _RAND_3505[7:0];
  _RAND_3506 = {1{`RANDOM}};
  lineBuffer_3499 = _RAND_3506[7:0];
  _RAND_3507 = {1{`RANDOM}};
  lineBuffer_3500 = _RAND_3507[7:0];
  _RAND_3508 = {1{`RANDOM}};
  lineBuffer_3501 = _RAND_3508[7:0];
  _RAND_3509 = {1{`RANDOM}};
  lineBuffer_3502 = _RAND_3509[7:0];
  _RAND_3510 = {1{`RANDOM}};
  lineBuffer_3503 = _RAND_3510[7:0];
  _RAND_3511 = {1{`RANDOM}};
  lineBuffer_3504 = _RAND_3511[7:0];
  _RAND_3512 = {1{`RANDOM}};
  lineBuffer_3505 = _RAND_3512[7:0];
  _RAND_3513 = {1{`RANDOM}};
  lineBuffer_3506 = _RAND_3513[7:0];
  _RAND_3514 = {1{`RANDOM}};
  lineBuffer_3507 = _RAND_3514[7:0];
  _RAND_3515 = {1{`RANDOM}};
  lineBuffer_3508 = _RAND_3515[7:0];
  _RAND_3516 = {1{`RANDOM}};
  lineBuffer_3509 = _RAND_3516[7:0];
  _RAND_3517 = {1{`RANDOM}};
  lineBuffer_3510 = _RAND_3517[7:0];
  _RAND_3518 = {1{`RANDOM}};
  lineBuffer_3511 = _RAND_3518[7:0];
  _RAND_3519 = {1{`RANDOM}};
  lineBuffer_3512 = _RAND_3519[7:0];
  _RAND_3520 = {1{`RANDOM}};
  lineBuffer_3513 = _RAND_3520[7:0];
  _RAND_3521 = {1{`RANDOM}};
  lineBuffer_3514 = _RAND_3521[7:0];
  _RAND_3522 = {1{`RANDOM}};
  lineBuffer_3515 = _RAND_3522[7:0];
  _RAND_3523 = {1{`RANDOM}};
  lineBuffer_3516 = _RAND_3523[7:0];
  _RAND_3524 = {1{`RANDOM}};
  lineBuffer_3517 = _RAND_3524[7:0];
  _RAND_3525 = {1{`RANDOM}};
  lineBuffer_3518 = _RAND_3525[7:0];
  _RAND_3526 = {1{`RANDOM}};
  lineBuffer_3519 = _RAND_3526[7:0];
  _RAND_3527 = {1{`RANDOM}};
  lineBuffer_3520 = _RAND_3527[7:0];
  _RAND_3528 = {1{`RANDOM}};
  lineBuffer_3521 = _RAND_3528[7:0];
  _RAND_3529 = {1{`RANDOM}};
  lineBuffer_3522 = _RAND_3529[7:0];
  _RAND_3530 = {1{`RANDOM}};
  lineBuffer_3523 = _RAND_3530[7:0];
  _RAND_3531 = {1{`RANDOM}};
  lineBuffer_3524 = _RAND_3531[7:0];
  _RAND_3532 = {1{`RANDOM}};
  lineBuffer_3525 = _RAND_3532[7:0];
  _RAND_3533 = {1{`RANDOM}};
  lineBuffer_3526 = _RAND_3533[7:0];
  _RAND_3534 = {1{`RANDOM}};
  lineBuffer_3527 = _RAND_3534[7:0];
  _RAND_3535 = {1{`RANDOM}};
  lineBuffer_3528 = _RAND_3535[7:0];
  _RAND_3536 = {1{`RANDOM}};
  lineBuffer_3529 = _RAND_3536[7:0];
  _RAND_3537 = {1{`RANDOM}};
  lineBuffer_3530 = _RAND_3537[7:0];
  _RAND_3538 = {1{`RANDOM}};
  lineBuffer_3531 = _RAND_3538[7:0];
  _RAND_3539 = {1{`RANDOM}};
  lineBuffer_3532 = _RAND_3539[7:0];
  _RAND_3540 = {1{`RANDOM}};
  lineBuffer_3533 = _RAND_3540[7:0];
  _RAND_3541 = {1{`RANDOM}};
  lineBuffer_3534 = _RAND_3541[7:0];
  _RAND_3542 = {1{`RANDOM}};
  lineBuffer_3535 = _RAND_3542[7:0];
  _RAND_3543 = {1{`RANDOM}};
  lineBuffer_3536 = _RAND_3543[7:0];
  _RAND_3544 = {1{`RANDOM}};
  lineBuffer_3537 = _RAND_3544[7:0];
  _RAND_3545 = {1{`RANDOM}};
  lineBuffer_3538 = _RAND_3545[7:0];
  _RAND_3546 = {1{`RANDOM}};
  lineBuffer_3539 = _RAND_3546[7:0];
  _RAND_3547 = {1{`RANDOM}};
  lineBuffer_3540 = _RAND_3547[7:0];
  _RAND_3548 = {1{`RANDOM}};
  lineBuffer_3541 = _RAND_3548[7:0];
  _RAND_3549 = {1{`RANDOM}};
  lineBuffer_3542 = _RAND_3549[7:0];
  _RAND_3550 = {1{`RANDOM}};
  lineBuffer_3543 = _RAND_3550[7:0];
  _RAND_3551 = {1{`RANDOM}};
  lineBuffer_3544 = _RAND_3551[7:0];
  _RAND_3552 = {1{`RANDOM}};
  lineBuffer_3545 = _RAND_3552[7:0];
  _RAND_3553 = {1{`RANDOM}};
  lineBuffer_3546 = _RAND_3553[7:0];
  _RAND_3554 = {1{`RANDOM}};
  lineBuffer_3547 = _RAND_3554[7:0];
  _RAND_3555 = {1{`RANDOM}};
  lineBuffer_3548 = _RAND_3555[7:0];
  _RAND_3556 = {1{`RANDOM}};
  lineBuffer_3549 = _RAND_3556[7:0];
  _RAND_3557 = {1{`RANDOM}};
  lineBuffer_3550 = _RAND_3557[7:0];
  _RAND_3558 = {1{`RANDOM}};
  lineBuffer_3551 = _RAND_3558[7:0];
  _RAND_3559 = {1{`RANDOM}};
  lineBuffer_3552 = _RAND_3559[7:0];
  _RAND_3560 = {1{`RANDOM}};
  lineBuffer_3553 = _RAND_3560[7:0];
  _RAND_3561 = {1{`RANDOM}};
  lineBuffer_3554 = _RAND_3561[7:0];
  _RAND_3562 = {1{`RANDOM}};
  lineBuffer_3555 = _RAND_3562[7:0];
  _RAND_3563 = {1{`RANDOM}};
  lineBuffer_3556 = _RAND_3563[7:0];
  _RAND_3564 = {1{`RANDOM}};
  lineBuffer_3557 = _RAND_3564[7:0];
  _RAND_3565 = {1{`RANDOM}};
  lineBuffer_3558 = _RAND_3565[7:0];
  _RAND_3566 = {1{`RANDOM}};
  lineBuffer_3559 = _RAND_3566[7:0];
  _RAND_3567 = {1{`RANDOM}};
  lineBuffer_3560 = _RAND_3567[7:0];
  _RAND_3568 = {1{`RANDOM}};
  lineBuffer_3561 = _RAND_3568[7:0];
  _RAND_3569 = {1{`RANDOM}};
  lineBuffer_3562 = _RAND_3569[7:0];
  _RAND_3570 = {1{`RANDOM}};
  lineBuffer_3563 = _RAND_3570[7:0];
  _RAND_3571 = {1{`RANDOM}};
  lineBuffer_3564 = _RAND_3571[7:0];
  _RAND_3572 = {1{`RANDOM}};
  lineBuffer_3565 = _RAND_3572[7:0];
  _RAND_3573 = {1{`RANDOM}};
  lineBuffer_3566 = _RAND_3573[7:0];
  _RAND_3574 = {1{`RANDOM}};
  lineBuffer_3567 = _RAND_3574[7:0];
  _RAND_3575 = {1{`RANDOM}};
  lineBuffer_3568 = _RAND_3575[7:0];
  _RAND_3576 = {1{`RANDOM}};
  lineBuffer_3569 = _RAND_3576[7:0];
  _RAND_3577 = {1{`RANDOM}};
  lineBuffer_3570 = _RAND_3577[7:0];
  _RAND_3578 = {1{`RANDOM}};
  lineBuffer_3571 = _RAND_3578[7:0];
  _RAND_3579 = {1{`RANDOM}};
  lineBuffer_3572 = _RAND_3579[7:0];
  _RAND_3580 = {1{`RANDOM}};
  lineBuffer_3573 = _RAND_3580[7:0];
  _RAND_3581 = {1{`RANDOM}};
  lineBuffer_3574 = _RAND_3581[7:0];
  _RAND_3582 = {1{`RANDOM}};
  lineBuffer_3575 = _RAND_3582[7:0];
  _RAND_3583 = {1{`RANDOM}};
  lineBuffer_3576 = _RAND_3583[7:0];
  _RAND_3584 = {1{`RANDOM}};
  lineBuffer_3577 = _RAND_3584[7:0];
  _RAND_3585 = {1{`RANDOM}};
  lineBuffer_3578 = _RAND_3585[7:0];
  _RAND_3586 = {1{`RANDOM}};
  lineBuffer_3579 = _RAND_3586[7:0];
  _RAND_3587 = {1{`RANDOM}};
  lineBuffer_3580 = _RAND_3587[7:0];
  _RAND_3588 = {1{`RANDOM}};
  lineBuffer_3581 = _RAND_3588[7:0];
  _RAND_3589 = {1{`RANDOM}};
  lineBuffer_3582 = _RAND_3589[7:0];
  _RAND_3590 = {1{`RANDOM}};
  lineBuffer_3583 = _RAND_3590[7:0];
  _RAND_3591 = {1{`RANDOM}};
  lineBuffer_3584 = _RAND_3591[7:0];
  _RAND_3592 = {1{`RANDOM}};
  lineBuffer_3585 = _RAND_3592[7:0];
  _RAND_3593 = {1{`RANDOM}};
  lineBuffer_3586 = _RAND_3593[7:0];
  _RAND_3594 = {1{`RANDOM}};
  lineBuffer_3587 = _RAND_3594[7:0];
  _RAND_3595 = {1{`RANDOM}};
  lineBuffer_3588 = _RAND_3595[7:0];
  _RAND_3596 = {1{`RANDOM}};
  lineBuffer_3589 = _RAND_3596[7:0];
  _RAND_3597 = {1{`RANDOM}};
  lineBuffer_3590 = _RAND_3597[7:0];
  _RAND_3598 = {1{`RANDOM}};
  lineBuffer_3591 = _RAND_3598[7:0];
  _RAND_3599 = {1{`RANDOM}};
  lineBuffer_3592 = _RAND_3599[7:0];
  _RAND_3600 = {1{`RANDOM}};
  lineBuffer_3593 = _RAND_3600[7:0];
  _RAND_3601 = {1{`RANDOM}};
  lineBuffer_3594 = _RAND_3601[7:0];
  _RAND_3602 = {1{`RANDOM}};
  lineBuffer_3595 = _RAND_3602[7:0];
  _RAND_3603 = {1{`RANDOM}};
  lineBuffer_3596 = _RAND_3603[7:0];
  _RAND_3604 = {1{`RANDOM}};
  lineBuffer_3597 = _RAND_3604[7:0];
  _RAND_3605 = {1{`RANDOM}};
  lineBuffer_3598 = _RAND_3605[7:0];
  _RAND_3606 = {1{`RANDOM}};
  lineBuffer_3599 = _RAND_3606[7:0];
  _RAND_3607 = {1{`RANDOM}};
  lineBuffer_3600 = _RAND_3607[7:0];
  _RAND_3608 = {1{`RANDOM}};
  lineBuffer_3601 = _RAND_3608[7:0];
  _RAND_3609 = {1{`RANDOM}};
  lineBuffer_3602 = _RAND_3609[7:0];
  _RAND_3610 = {1{`RANDOM}};
  lineBuffer_3603 = _RAND_3610[7:0];
  _RAND_3611 = {1{`RANDOM}};
  lineBuffer_3604 = _RAND_3611[7:0];
  _RAND_3612 = {1{`RANDOM}};
  lineBuffer_3605 = _RAND_3612[7:0];
  _RAND_3613 = {1{`RANDOM}};
  lineBuffer_3606 = _RAND_3613[7:0];
  _RAND_3614 = {1{`RANDOM}};
  lineBuffer_3607 = _RAND_3614[7:0];
  _RAND_3615 = {1{`RANDOM}};
  lineBuffer_3608 = _RAND_3615[7:0];
  _RAND_3616 = {1{`RANDOM}};
  lineBuffer_3609 = _RAND_3616[7:0];
  _RAND_3617 = {1{`RANDOM}};
  lineBuffer_3610 = _RAND_3617[7:0];
  _RAND_3618 = {1{`RANDOM}};
  lineBuffer_3611 = _RAND_3618[7:0];
  _RAND_3619 = {1{`RANDOM}};
  lineBuffer_3612 = _RAND_3619[7:0];
  _RAND_3620 = {1{`RANDOM}};
  lineBuffer_3613 = _RAND_3620[7:0];
  _RAND_3621 = {1{`RANDOM}};
  lineBuffer_3614 = _RAND_3621[7:0];
  _RAND_3622 = {1{`RANDOM}};
  lineBuffer_3615 = _RAND_3622[7:0];
  _RAND_3623 = {1{`RANDOM}};
  lineBuffer_3616 = _RAND_3623[7:0];
  _RAND_3624 = {1{`RANDOM}};
  lineBuffer_3617 = _RAND_3624[7:0];
  _RAND_3625 = {1{`RANDOM}};
  lineBuffer_3618 = _RAND_3625[7:0];
  _RAND_3626 = {1{`RANDOM}};
  lineBuffer_3619 = _RAND_3626[7:0];
  _RAND_3627 = {1{`RANDOM}};
  lineBuffer_3620 = _RAND_3627[7:0];
  _RAND_3628 = {1{`RANDOM}};
  lineBuffer_3621 = _RAND_3628[7:0];
  _RAND_3629 = {1{`RANDOM}};
  lineBuffer_3622 = _RAND_3629[7:0];
  _RAND_3630 = {1{`RANDOM}};
  lineBuffer_3623 = _RAND_3630[7:0];
  _RAND_3631 = {1{`RANDOM}};
  lineBuffer_3624 = _RAND_3631[7:0];
  _RAND_3632 = {1{`RANDOM}};
  lineBuffer_3625 = _RAND_3632[7:0];
  _RAND_3633 = {1{`RANDOM}};
  lineBuffer_3626 = _RAND_3633[7:0];
  _RAND_3634 = {1{`RANDOM}};
  lineBuffer_3627 = _RAND_3634[7:0];
  _RAND_3635 = {1{`RANDOM}};
  lineBuffer_3628 = _RAND_3635[7:0];
  _RAND_3636 = {1{`RANDOM}};
  lineBuffer_3629 = _RAND_3636[7:0];
  _RAND_3637 = {1{`RANDOM}};
  lineBuffer_3630 = _RAND_3637[7:0];
  _RAND_3638 = {1{`RANDOM}};
  lineBuffer_3631 = _RAND_3638[7:0];
  _RAND_3639 = {1{`RANDOM}};
  lineBuffer_3632 = _RAND_3639[7:0];
  _RAND_3640 = {1{`RANDOM}};
  lineBuffer_3633 = _RAND_3640[7:0];
  _RAND_3641 = {1{`RANDOM}};
  lineBuffer_3634 = _RAND_3641[7:0];
  _RAND_3642 = {1{`RANDOM}};
  lineBuffer_3635 = _RAND_3642[7:0];
  _RAND_3643 = {1{`RANDOM}};
  lineBuffer_3636 = _RAND_3643[7:0];
  _RAND_3644 = {1{`RANDOM}};
  lineBuffer_3637 = _RAND_3644[7:0];
  _RAND_3645 = {1{`RANDOM}};
  lineBuffer_3638 = _RAND_3645[7:0];
  _RAND_3646 = {1{`RANDOM}};
  lineBuffer_3639 = _RAND_3646[7:0];
  _RAND_3647 = {1{`RANDOM}};
  lineBuffer_3640 = _RAND_3647[7:0];
  _RAND_3648 = {1{`RANDOM}};
  lineBuffer_3641 = _RAND_3648[7:0];
  _RAND_3649 = {1{`RANDOM}};
  lineBuffer_3642 = _RAND_3649[7:0];
  _RAND_3650 = {1{`RANDOM}};
  lineBuffer_3643 = _RAND_3650[7:0];
  _RAND_3651 = {1{`RANDOM}};
  lineBuffer_3644 = _RAND_3651[7:0];
  _RAND_3652 = {1{`RANDOM}};
  lineBuffer_3645 = _RAND_3652[7:0];
  _RAND_3653 = {1{`RANDOM}};
  lineBuffer_3646 = _RAND_3653[7:0];
  _RAND_3654 = {1{`RANDOM}};
  lineBuffer_3647 = _RAND_3654[7:0];
  _RAND_3655 = {1{`RANDOM}};
  lineBuffer_3648 = _RAND_3655[7:0];
  _RAND_3656 = {1{`RANDOM}};
  lineBuffer_3649 = _RAND_3656[7:0];
  _RAND_3657 = {1{`RANDOM}};
  lineBuffer_3650 = _RAND_3657[7:0];
  _RAND_3658 = {1{`RANDOM}};
  lineBuffer_3651 = _RAND_3658[7:0];
  _RAND_3659 = {1{`RANDOM}};
  lineBuffer_3652 = _RAND_3659[7:0];
  _RAND_3660 = {1{`RANDOM}};
  lineBuffer_3653 = _RAND_3660[7:0];
  _RAND_3661 = {1{`RANDOM}};
  lineBuffer_3654 = _RAND_3661[7:0];
  _RAND_3662 = {1{`RANDOM}};
  lineBuffer_3655 = _RAND_3662[7:0];
  _RAND_3663 = {1{`RANDOM}};
  lineBuffer_3656 = _RAND_3663[7:0];
  _RAND_3664 = {1{`RANDOM}};
  lineBuffer_3657 = _RAND_3664[7:0];
  _RAND_3665 = {1{`RANDOM}};
  lineBuffer_3658 = _RAND_3665[7:0];
  _RAND_3666 = {1{`RANDOM}};
  lineBuffer_3659 = _RAND_3666[7:0];
  _RAND_3667 = {1{`RANDOM}};
  lineBuffer_3660 = _RAND_3667[7:0];
  _RAND_3668 = {1{`RANDOM}};
  lineBuffer_3661 = _RAND_3668[7:0];
  _RAND_3669 = {1{`RANDOM}};
  lineBuffer_3662 = _RAND_3669[7:0];
  _RAND_3670 = {1{`RANDOM}};
  lineBuffer_3663 = _RAND_3670[7:0];
  _RAND_3671 = {1{`RANDOM}};
  lineBuffer_3664 = _RAND_3671[7:0];
  _RAND_3672 = {1{`RANDOM}};
  lineBuffer_3665 = _RAND_3672[7:0];
  _RAND_3673 = {1{`RANDOM}};
  lineBuffer_3666 = _RAND_3673[7:0];
  _RAND_3674 = {1{`RANDOM}};
  lineBuffer_3667 = _RAND_3674[7:0];
  _RAND_3675 = {1{`RANDOM}};
  lineBuffer_3668 = _RAND_3675[7:0];
  _RAND_3676 = {1{`RANDOM}};
  lineBuffer_3669 = _RAND_3676[7:0];
  _RAND_3677 = {1{`RANDOM}};
  lineBuffer_3670 = _RAND_3677[7:0];
  _RAND_3678 = {1{`RANDOM}};
  lineBuffer_3671 = _RAND_3678[7:0];
  _RAND_3679 = {1{`RANDOM}};
  lineBuffer_3672 = _RAND_3679[7:0];
  _RAND_3680 = {1{`RANDOM}};
  lineBuffer_3673 = _RAND_3680[7:0];
  _RAND_3681 = {1{`RANDOM}};
  lineBuffer_3674 = _RAND_3681[7:0];
  _RAND_3682 = {1{`RANDOM}};
  lineBuffer_3675 = _RAND_3682[7:0];
  _RAND_3683 = {1{`RANDOM}};
  lineBuffer_3676 = _RAND_3683[7:0];
  _RAND_3684 = {1{`RANDOM}};
  lineBuffer_3677 = _RAND_3684[7:0];
  _RAND_3685 = {1{`RANDOM}};
  lineBuffer_3678 = _RAND_3685[7:0];
  _RAND_3686 = {1{`RANDOM}};
  lineBuffer_3679 = _RAND_3686[7:0];
  _RAND_3687 = {1{`RANDOM}};
  lineBuffer_3680 = _RAND_3687[7:0];
  _RAND_3688 = {1{`RANDOM}};
  lineBuffer_3681 = _RAND_3688[7:0];
  _RAND_3689 = {1{`RANDOM}};
  lineBuffer_3682 = _RAND_3689[7:0];
  _RAND_3690 = {1{`RANDOM}};
  lineBuffer_3683 = _RAND_3690[7:0];
  _RAND_3691 = {1{`RANDOM}};
  lineBuffer_3684 = _RAND_3691[7:0];
  _RAND_3692 = {1{`RANDOM}};
  lineBuffer_3685 = _RAND_3692[7:0];
  _RAND_3693 = {1{`RANDOM}};
  lineBuffer_3686 = _RAND_3693[7:0];
  _RAND_3694 = {1{`RANDOM}};
  lineBuffer_3687 = _RAND_3694[7:0];
  _RAND_3695 = {1{`RANDOM}};
  lineBuffer_3688 = _RAND_3695[7:0];
  _RAND_3696 = {1{`RANDOM}};
  lineBuffer_3689 = _RAND_3696[7:0];
  _RAND_3697 = {1{`RANDOM}};
  lineBuffer_3690 = _RAND_3697[7:0];
  _RAND_3698 = {1{`RANDOM}};
  lineBuffer_3691 = _RAND_3698[7:0];
  _RAND_3699 = {1{`RANDOM}};
  lineBuffer_3692 = _RAND_3699[7:0];
  _RAND_3700 = {1{`RANDOM}};
  lineBuffer_3693 = _RAND_3700[7:0];
  _RAND_3701 = {1{`RANDOM}};
  lineBuffer_3694 = _RAND_3701[7:0];
  _RAND_3702 = {1{`RANDOM}};
  lineBuffer_3695 = _RAND_3702[7:0];
  _RAND_3703 = {1{`RANDOM}};
  lineBuffer_3696 = _RAND_3703[7:0];
  _RAND_3704 = {1{`RANDOM}};
  lineBuffer_3697 = _RAND_3704[7:0];
  _RAND_3705 = {1{`RANDOM}};
  lineBuffer_3698 = _RAND_3705[7:0];
  _RAND_3706 = {1{`RANDOM}};
  lineBuffer_3699 = _RAND_3706[7:0];
  _RAND_3707 = {1{`RANDOM}};
  lineBuffer_3700 = _RAND_3707[7:0];
  _RAND_3708 = {1{`RANDOM}};
  lineBuffer_3701 = _RAND_3708[7:0];
  _RAND_3709 = {1{`RANDOM}};
  lineBuffer_3702 = _RAND_3709[7:0];
  _RAND_3710 = {1{`RANDOM}};
  lineBuffer_3703 = _RAND_3710[7:0];
  _RAND_3711 = {1{`RANDOM}};
  lineBuffer_3704 = _RAND_3711[7:0];
  _RAND_3712 = {1{`RANDOM}};
  lineBuffer_3705 = _RAND_3712[7:0];
  _RAND_3713 = {1{`RANDOM}};
  lineBuffer_3706 = _RAND_3713[7:0];
  _RAND_3714 = {1{`RANDOM}};
  lineBuffer_3707 = _RAND_3714[7:0];
  _RAND_3715 = {1{`RANDOM}};
  lineBuffer_3708 = _RAND_3715[7:0];
  _RAND_3716 = {1{`RANDOM}};
  lineBuffer_3709 = _RAND_3716[7:0];
  _RAND_3717 = {1{`RANDOM}};
  lineBuffer_3710 = _RAND_3717[7:0];
  _RAND_3718 = {1{`RANDOM}};
  lineBuffer_3711 = _RAND_3718[7:0];
  _RAND_3719 = {1{`RANDOM}};
  lineBuffer_3712 = _RAND_3719[7:0];
  _RAND_3720 = {1{`RANDOM}};
  lineBuffer_3713 = _RAND_3720[7:0];
  _RAND_3721 = {1{`RANDOM}};
  lineBuffer_3714 = _RAND_3721[7:0];
  _RAND_3722 = {1{`RANDOM}};
  lineBuffer_3715 = _RAND_3722[7:0];
  _RAND_3723 = {1{`RANDOM}};
  lineBuffer_3716 = _RAND_3723[7:0];
  _RAND_3724 = {1{`RANDOM}};
  lineBuffer_3717 = _RAND_3724[7:0];
  _RAND_3725 = {1{`RANDOM}};
  lineBuffer_3718 = _RAND_3725[7:0];
  _RAND_3726 = {1{`RANDOM}};
  lineBuffer_3719 = _RAND_3726[7:0];
  _RAND_3727 = {1{`RANDOM}};
  lineBuffer_3720 = _RAND_3727[7:0];
  _RAND_3728 = {1{`RANDOM}};
  lineBuffer_3721 = _RAND_3728[7:0];
  _RAND_3729 = {1{`RANDOM}};
  lineBuffer_3722 = _RAND_3729[7:0];
  _RAND_3730 = {1{`RANDOM}};
  lineBuffer_3723 = _RAND_3730[7:0];
  _RAND_3731 = {1{`RANDOM}};
  lineBuffer_3724 = _RAND_3731[7:0];
  _RAND_3732 = {1{`RANDOM}};
  lineBuffer_3725 = _RAND_3732[7:0];
  _RAND_3733 = {1{`RANDOM}};
  lineBuffer_3726 = _RAND_3733[7:0];
  _RAND_3734 = {1{`RANDOM}};
  lineBuffer_3727 = _RAND_3734[7:0];
  _RAND_3735 = {1{`RANDOM}};
  lineBuffer_3728 = _RAND_3735[7:0];
  _RAND_3736 = {1{`RANDOM}};
  lineBuffer_3729 = _RAND_3736[7:0];
  _RAND_3737 = {1{`RANDOM}};
  lineBuffer_3730 = _RAND_3737[7:0];
  _RAND_3738 = {1{`RANDOM}};
  lineBuffer_3731 = _RAND_3738[7:0];
  _RAND_3739 = {1{`RANDOM}};
  lineBuffer_3732 = _RAND_3739[7:0];
  _RAND_3740 = {1{`RANDOM}};
  lineBuffer_3733 = _RAND_3740[7:0];
  _RAND_3741 = {1{`RANDOM}};
  lineBuffer_3734 = _RAND_3741[7:0];
  _RAND_3742 = {1{`RANDOM}};
  lineBuffer_3735 = _RAND_3742[7:0];
  _RAND_3743 = {1{`RANDOM}};
  lineBuffer_3736 = _RAND_3743[7:0];
  _RAND_3744 = {1{`RANDOM}};
  lineBuffer_3737 = _RAND_3744[7:0];
  _RAND_3745 = {1{`RANDOM}};
  lineBuffer_3738 = _RAND_3745[7:0];
  _RAND_3746 = {1{`RANDOM}};
  lineBuffer_3739 = _RAND_3746[7:0];
  _RAND_3747 = {1{`RANDOM}};
  lineBuffer_3740 = _RAND_3747[7:0];
  _RAND_3748 = {1{`RANDOM}};
  lineBuffer_3741 = _RAND_3748[7:0];
  _RAND_3749 = {1{`RANDOM}};
  lineBuffer_3742 = _RAND_3749[7:0];
  _RAND_3750 = {1{`RANDOM}};
  lineBuffer_3743 = _RAND_3750[7:0];
  _RAND_3751 = {1{`RANDOM}};
  lineBuffer_3744 = _RAND_3751[7:0];
  _RAND_3752 = {1{`RANDOM}};
  lineBuffer_3745 = _RAND_3752[7:0];
  _RAND_3753 = {1{`RANDOM}};
  lineBuffer_3746 = _RAND_3753[7:0];
  _RAND_3754 = {1{`RANDOM}};
  lineBuffer_3747 = _RAND_3754[7:0];
  _RAND_3755 = {1{`RANDOM}};
  lineBuffer_3748 = _RAND_3755[7:0];
  _RAND_3756 = {1{`RANDOM}};
  lineBuffer_3749 = _RAND_3756[7:0];
  _RAND_3757 = {1{`RANDOM}};
  lineBuffer_3750 = _RAND_3757[7:0];
  _RAND_3758 = {1{`RANDOM}};
  lineBuffer_3751 = _RAND_3758[7:0];
  _RAND_3759 = {1{`RANDOM}};
  lineBuffer_3752 = _RAND_3759[7:0];
  _RAND_3760 = {1{`RANDOM}};
  lineBuffer_3753 = _RAND_3760[7:0];
  _RAND_3761 = {1{`RANDOM}};
  lineBuffer_3754 = _RAND_3761[7:0];
  _RAND_3762 = {1{`RANDOM}};
  lineBuffer_3755 = _RAND_3762[7:0];
  _RAND_3763 = {1{`RANDOM}};
  lineBuffer_3756 = _RAND_3763[7:0];
  _RAND_3764 = {1{`RANDOM}};
  lineBuffer_3757 = _RAND_3764[7:0];
  _RAND_3765 = {1{`RANDOM}};
  lineBuffer_3758 = _RAND_3765[7:0];
  _RAND_3766 = {1{`RANDOM}};
  lineBuffer_3759 = _RAND_3766[7:0];
  _RAND_3767 = {1{`RANDOM}};
  lineBuffer_3760 = _RAND_3767[7:0];
  _RAND_3768 = {1{`RANDOM}};
  lineBuffer_3761 = _RAND_3768[7:0];
  _RAND_3769 = {1{`RANDOM}};
  lineBuffer_3762 = _RAND_3769[7:0];
  _RAND_3770 = {1{`RANDOM}};
  lineBuffer_3763 = _RAND_3770[7:0];
  _RAND_3771 = {1{`RANDOM}};
  lineBuffer_3764 = _RAND_3771[7:0];
  _RAND_3772 = {1{`RANDOM}};
  lineBuffer_3765 = _RAND_3772[7:0];
  _RAND_3773 = {1{`RANDOM}};
  lineBuffer_3766 = _RAND_3773[7:0];
  _RAND_3774 = {1{`RANDOM}};
  lineBuffer_3767 = _RAND_3774[7:0];
  _RAND_3775 = {1{`RANDOM}};
  lineBuffer_3768 = _RAND_3775[7:0];
  _RAND_3776 = {1{`RANDOM}};
  lineBuffer_3769 = _RAND_3776[7:0];
  _RAND_3777 = {1{`RANDOM}};
  lineBuffer_3770 = _RAND_3777[7:0];
  _RAND_3778 = {1{`RANDOM}};
  lineBuffer_3771 = _RAND_3778[7:0];
  _RAND_3779 = {1{`RANDOM}};
  lineBuffer_3772 = _RAND_3779[7:0];
  _RAND_3780 = {1{`RANDOM}};
  lineBuffer_3773 = _RAND_3780[7:0];
  _RAND_3781 = {1{`RANDOM}};
  lineBuffer_3774 = _RAND_3781[7:0];
  _RAND_3782 = {1{`RANDOM}};
  lineBuffer_3775 = _RAND_3782[7:0];
  _RAND_3783 = {1{`RANDOM}};
  lineBuffer_3776 = _RAND_3783[7:0];
  _RAND_3784 = {1{`RANDOM}};
  lineBuffer_3777 = _RAND_3784[7:0];
  _RAND_3785 = {1{`RANDOM}};
  lineBuffer_3778 = _RAND_3785[7:0];
  _RAND_3786 = {1{`RANDOM}};
  lineBuffer_3779 = _RAND_3786[7:0];
  _RAND_3787 = {1{`RANDOM}};
  lineBuffer_3780 = _RAND_3787[7:0];
  _RAND_3788 = {1{`RANDOM}};
  lineBuffer_3781 = _RAND_3788[7:0];
  _RAND_3789 = {1{`RANDOM}};
  lineBuffer_3782 = _RAND_3789[7:0];
  _RAND_3790 = {1{`RANDOM}};
  lineBuffer_3783 = _RAND_3790[7:0];
  _RAND_3791 = {1{`RANDOM}};
  lineBuffer_3784 = _RAND_3791[7:0];
  _RAND_3792 = {1{`RANDOM}};
  lineBuffer_3785 = _RAND_3792[7:0];
  _RAND_3793 = {1{`RANDOM}};
  lineBuffer_3786 = _RAND_3793[7:0];
  _RAND_3794 = {1{`RANDOM}};
  lineBuffer_3787 = _RAND_3794[7:0];
  _RAND_3795 = {1{`RANDOM}};
  lineBuffer_3788 = _RAND_3795[7:0];
  _RAND_3796 = {1{`RANDOM}};
  lineBuffer_3789 = _RAND_3796[7:0];
  _RAND_3797 = {1{`RANDOM}};
  lineBuffer_3790 = _RAND_3797[7:0];
  _RAND_3798 = {1{`RANDOM}};
  lineBuffer_3791 = _RAND_3798[7:0];
  _RAND_3799 = {1{`RANDOM}};
  lineBuffer_3792 = _RAND_3799[7:0];
  _RAND_3800 = {1{`RANDOM}};
  lineBuffer_3793 = _RAND_3800[7:0];
  _RAND_3801 = {1{`RANDOM}};
  lineBuffer_3794 = _RAND_3801[7:0];
  _RAND_3802 = {1{`RANDOM}};
  lineBuffer_3795 = _RAND_3802[7:0];
  _RAND_3803 = {1{`RANDOM}};
  lineBuffer_3796 = _RAND_3803[7:0];
  _RAND_3804 = {1{`RANDOM}};
  lineBuffer_3797 = _RAND_3804[7:0];
  _RAND_3805 = {1{`RANDOM}};
  lineBuffer_3798 = _RAND_3805[7:0];
  _RAND_3806 = {1{`RANDOM}};
  lineBuffer_3799 = _RAND_3806[7:0];
  _RAND_3807 = {1{`RANDOM}};
  lineBuffer_3800 = _RAND_3807[7:0];
  _RAND_3808 = {1{`RANDOM}};
  lineBuffer_3801 = _RAND_3808[7:0];
  _RAND_3809 = {1{`RANDOM}};
  lineBuffer_3802 = _RAND_3809[7:0];
  _RAND_3810 = {1{`RANDOM}};
  lineBuffer_3803 = _RAND_3810[7:0];
  _RAND_3811 = {1{`RANDOM}};
  lineBuffer_3804 = _RAND_3811[7:0];
  _RAND_3812 = {1{`RANDOM}};
  lineBuffer_3805 = _RAND_3812[7:0];
  _RAND_3813 = {1{`RANDOM}};
  lineBuffer_3806 = _RAND_3813[7:0];
  _RAND_3814 = {1{`RANDOM}};
  lineBuffer_3807 = _RAND_3814[7:0];
  _RAND_3815 = {1{`RANDOM}};
  lineBuffer_3808 = _RAND_3815[7:0];
  _RAND_3816 = {1{`RANDOM}};
  lineBuffer_3809 = _RAND_3816[7:0];
  _RAND_3817 = {1{`RANDOM}};
  lineBuffer_3810 = _RAND_3817[7:0];
  _RAND_3818 = {1{`RANDOM}};
  lineBuffer_3811 = _RAND_3818[7:0];
  _RAND_3819 = {1{`RANDOM}};
  lineBuffer_3812 = _RAND_3819[7:0];
  _RAND_3820 = {1{`RANDOM}};
  lineBuffer_3813 = _RAND_3820[7:0];
  _RAND_3821 = {1{`RANDOM}};
  lineBuffer_3814 = _RAND_3821[7:0];
  _RAND_3822 = {1{`RANDOM}};
  lineBuffer_3815 = _RAND_3822[7:0];
  _RAND_3823 = {1{`RANDOM}};
  lineBuffer_3816 = _RAND_3823[7:0];
  _RAND_3824 = {1{`RANDOM}};
  lineBuffer_3817 = _RAND_3824[7:0];
  _RAND_3825 = {1{`RANDOM}};
  lineBuffer_3818 = _RAND_3825[7:0];
  _RAND_3826 = {1{`RANDOM}};
  lineBuffer_3819 = _RAND_3826[7:0];
  _RAND_3827 = {1{`RANDOM}};
  lineBuffer_3820 = _RAND_3827[7:0];
  _RAND_3828 = {1{`RANDOM}};
  lineBuffer_3821 = _RAND_3828[7:0];
  _RAND_3829 = {1{`RANDOM}};
  lineBuffer_3822 = _RAND_3829[7:0];
  _RAND_3830 = {1{`RANDOM}};
  lineBuffer_3823 = _RAND_3830[7:0];
  _RAND_3831 = {1{`RANDOM}};
  lineBuffer_3824 = _RAND_3831[7:0];
  _RAND_3832 = {1{`RANDOM}};
  lineBuffer_3825 = _RAND_3832[7:0];
  _RAND_3833 = {1{`RANDOM}};
  lineBuffer_3826 = _RAND_3833[7:0];
  _RAND_3834 = {1{`RANDOM}};
  lineBuffer_3827 = _RAND_3834[7:0];
  _RAND_3835 = {1{`RANDOM}};
  lineBuffer_3828 = _RAND_3835[7:0];
  _RAND_3836 = {1{`RANDOM}};
  lineBuffer_3829 = _RAND_3836[7:0];
  _RAND_3837 = {1{`RANDOM}};
  lineBuffer_3830 = _RAND_3837[7:0];
  _RAND_3838 = {1{`RANDOM}};
  lineBuffer_3831 = _RAND_3838[7:0];
  _RAND_3839 = {1{`RANDOM}};
  lineBuffer_3832 = _RAND_3839[7:0];
  _RAND_3840 = {1{`RANDOM}};
  lineBuffer_3833 = _RAND_3840[7:0];
  _RAND_3841 = {1{`RANDOM}};
  lineBuffer_3834 = _RAND_3841[7:0];
  _RAND_3842 = {1{`RANDOM}};
  lineBuffer_3835 = _RAND_3842[7:0];
  _RAND_3843 = {1{`RANDOM}};
  lineBuffer_3836 = _RAND_3843[7:0];
  _RAND_3844 = {1{`RANDOM}};
  lineBuffer_3837 = _RAND_3844[7:0];
  _RAND_3845 = {1{`RANDOM}};
  lineBuffer_3838 = _RAND_3845[7:0];
  _RAND_3846 = {1{`RANDOM}};
  lineBuffer_3839 = _RAND_3846[7:0];
  _RAND_3847 = {1{`RANDOM}};
  lineBuffer_3840 = _RAND_3847[7:0];
  _RAND_3848 = {1{`RANDOM}};
  lineBuffer_3841 = _RAND_3848[7:0];
  _RAND_3849 = {1{`RANDOM}};
  lineBuffer_3842 = _RAND_3849[7:0];
  _RAND_3850 = {1{`RANDOM}};
  lineBuffer_3843 = _RAND_3850[7:0];
  _RAND_3851 = {1{`RANDOM}};
  lineBuffer_3844 = _RAND_3851[7:0];
  _RAND_3852 = {1{`RANDOM}};
  lineBuffer_3845 = _RAND_3852[7:0];
  _RAND_3853 = {1{`RANDOM}};
  lineBuffer_3846 = _RAND_3853[7:0];
  _RAND_3854 = {1{`RANDOM}};
  lineBuffer_3847 = _RAND_3854[7:0];
  _RAND_3855 = {1{`RANDOM}};
  lineBuffer_3848 = _RAND_3855[7:0];
  _RAND_3856 = {1{`RANDOM}};
  lineBuffer_3849 = _RAND_3856[7:0];
  _RAND_3857 = {1{`RANDOM}};
  lineBuffer_3850 = _RAND_3857[7:0];
  _RAND_3858 = {1{`RANDOM}};
  lineBuffer_3851 = _RAND_3858[7:0];
  _RAND_3859 = {1{`RANDOM}};
  lineBuffer_3852 = _RAND_3859[7:0];
  _RAND_3860 = {1{`RANDOM}};
  lineBuffer_3853 = _RAND_3860[7:0];
  _RAND_3861 = {1{`RANDOM}};
  lineBuffer_3854 = _RAND_3861[7:0];
  _RAND_3862 = {1{`RANDOM}};
  lineBuffer_3855 = _RAND_3862[7:0];
  _RAND_3863 = {1{`RANDOM}};
  lineBuffer_3856 = _RAND_3863[7:0];
  _RAND_3864 = {1{`RANDOM}};
  lineBuffer_3857 = _RAND_3864[7:0];
  _RAND_3865 = {1{`RANDOM}};
  lineBuffer_3858 = _RAND_3865[7:0];
  _RAND_3866 = {1{`RANDOM}};
  lineBuffer_3859 = _RAND_3866[7:0];
  _RAND_3867 = {1{`RANDOM}};
  lineBuffer_3860 = _RAND_3867[7:0];
  _RAND_3868 = {1{`RANDOM}};
  lineBuffer_3861 = _RAND_3868[7:0];
  _RAND_3869 = {1{`RANDOM}};
  lineBuffer_3862 = _RAND_3869[7:0];
  _RAND_3870 = {1{`RANDOM}};
  lineBuffer_3863 = _RAND_3870[7:0];
  _RAND_3871 = {1{`RANDOM}};
  lineBuffer_3864 = _RAND_3871[7:0];
  _RAND_3872 = {1{`RANDOM}};
  lineBuffer_3865 = _RAND_3872[7:0];
  _RAND_3873 = {1{`RANDOM}};
  lineBuffer_3866 = _RAND_3873[7:0];
  _RAND_3874 = {1{`RANDOM}};
  lineBuffer_3867 = _RAND_3874[7:0];
  _RAND_3875 = {1{`RANDOM}};
  lineBuffer_3868 = _RAND_3875[7:0];
  _RAND_3876 = {1{`RANDOM}};
  lineBuffer_3869 = _RAND_3876[7:0];
  _RAND_3877 = {1{`RANDOM}};
  lineBuffer_3870 = _RAND_3877[7:0];
  _RAND_3878 = {1{`RANDOM}};
  lineBuffer_3871 = _RAND_3878[7:0];
  _RAND_3879 = {1{`RANDOM}};
  lineBuffer_3872 = _RAND_3879[7:0];
  _RAND_3880 = {1{`RANDOM}};
  lineBuffer_3873 = _RAND_3880[7:0];
  _RAND_3881 = {1{`RANDOM}};
  lineBuffer_3874 = _RAND_3881[7:0];
  _RAND_3882 = {1{`RANDOM}};
  lineBuffer_3875 = _RAND_3882[7:0];
  _RAND_3883 = {1{`RANDOM}};
  lineBuffer_3876 = _RAND_3883[7:0];
  _RAND_3884 = {1{`RANDOM}};
  lineBuffer_3877 = _RAND_3884[7:0];
  _RAND_3885 = {1{`RANDOM}};
  lineBuffer_3878 = _RAND_3885[7:0];
  _RAND_3886 = {1{`RANDOM}};
  lineBuffer_3879 = _RAND_3886[7:0];
  _RAND_3887 = {1{`RANDOM}};
  lineBuffer_3880 = _RAND_3887[7:0];
  _RAND_3888 = {1{`RANDOM}};
  lineBuffer_3881 = _RAND_3888[7:0];
  _RAND_3889 = {1{`RANDOM}};
  lineBuffer_3882 = _RAND_3889[7:0];
  _RAND_3890 = {1{`RANDOM}};
  lineBuffer_3883 = _RAND_3890[7:0];
  _RAND_3891 = {1{`RANDOM}};
  lineBuffer_3884 = _RAND_3891[7:0];
  _RAND_3892 = {1{`RANDOM}};
  lineBuffer_3885 = _RAND_3892[7:0];
  _RAND_3893 = {1{`RANDOM}};
  lineBuffer_3886 = _RAND_3893[7:0];
  _RAND_3894 = {1{`RANDOM}};
  lineBuffer_3887 = _RAND_3894[7:0];
  _RAND_3895 = {1{`RANDOM}};
  lineBuffer_3888 = _RAND_3895[7:0];
  _RAND_3896 = {1{`RANDOM}};
  lineBuffer_3889 = _RAND_3896[7:0];
  _RAND_3897 = {1{`RANDOM}};
  lineBuffer_3890 = _RAND_3897[7:0];
  _RAND_3898 = {1{`RANDOM}};
  lineBuffer_3891 = _RAND_3898[7:0];
  _RAND_3899 = {1{`RANDOM}};
  lineBuffer_3892 = _RAND_3899[7:0];
  _RAND_3900 = {1{`RANDOM}};
  lineBuffer_3893 = _RAND_3900[7:0];
  _RAND_3901 = {1{`RANDOM}};
  lineBuffer_3894 = _RAND_3901[7:0];
  _RAND_3902 = {1{`RANDOM}};
  lineBuffer_3895 = _RAND_3902[7:0];
  _RAND_3903 = {1{`RANDOM}};
  lineBuffer_3896 = _RAND_3903[7:0];
  _RAND_3904 = {1{`RANDOM}};
  lineBuffer_3897 = _RAND_3904[7:0];
  _RAND_3905 = {1{`RANDOM}};
  lineBuffer_3898 = _RAND_3905[7:0];
  _RAND_3906 = {1{`RANDOM}};
  lineBuffer_3899 = _RAND_3906[7:0];
  _RAND_3907 = {1{`RANDOM}};
  lineBuffer_3900 = _RAND_3907[7:0];
  _RAND_3908 = {1{`RANDOM}};
  lineBuffer_3901 = _RAND_3908[7:0];
  _RAND_3909 = {1{`RANDOM}};
  lineBuffer_3902 = _RAND_3909[7:0];
  _RAND_3910 = {1{`RANDOM}};
  lineBuffer_3903 = _RAND_3910[7:0];
  _RAND_3911 = {1{`RANDOM}};
  lineBuffer_3904 = _RAND_3911[7:0];
  _RAND_3912 = {1{`RANDOM}};
  lineBuffer_3905 = _RAND_3912[7:0];
  _RAND_3913 = {1{`RANDOM}};
  lineBuffer_3906 = _RAND_3913[7:0];
  _RAND_3914 = {1{`RANDOM}};
  lineBuffer_3907 = _RAND_3914[7:0];
  _RAND_3915 = {1{`RANDOM}};
  lineBuffer_3908 = _RAND_3915[7:0];
  _RAND_3916 = {1{`RANDOM}};
  lineBuffer_3909 = _RAND_3916[7:0];
  _RAND_3917 = {1{`RANDOM}};
  lineBuffer_3910 = _RAND_3917[7:0];
  _RAND_3918 = {1{`RANDOM}};
  lineBuffer_3911 = _RAND_3918[7:0];
  _RAND_3919 = {1{`RANDOM}};
  lineBuffer_3912 = _RAND_3919[7:0];
  _RAND_3920 = {1{`RANDOM}};
  lineBuffer_3913 = _RAND_3920[7:0];
  _RAND_3921 = {1{`RANDOM}};
  lineBuffer_3914 = _RAND_3921[7:0];
  _RAND_3922 = {1{`RANDOM}};
  lineBuffer_3915 = _RAND_3922[7:0];
  _RAND_3923 = {1{`RANDOM}};
  lineBuffer_3916 = _RAND_3923[7:0];
  _RAND_3924 = {1{`RANDOM}};
  lineBuffer_3917 = _RAND_3924[7:0];
  _RAND_3925 = {1{`RANDOM}};
  lineBuffer_3918 = _RAND_3925[7:0];
  _RAND_3926 = {1{`RANDOM}};
  lineBuffer_3919 = _RAND_3926[7:0];
  _RAND_3927 = {1{`RANDOM}};
  lineBuffer_3920 = _RAND_3927[7:0];
  _RAND_3928 = {1{`RANDOM}};
  lineBuffer_3921 = _RAND_3928[7:0];
  _RAND_3929 = {1{`RANDOM}};
  lineBuffer_3922 = _RAND_3929[7:0];
  _RAND_3930 = {1{`RANDOM}};
  lineBuffer_3923 = _RAND_3930[7:0];
  _RAND_3931 = {1{`RANDOM}};
  lineBuffer_3924 = _RAND_3931[7:0];
  _RAND_3932 = {1{`RANDOM}};
  lineBuffer_3925 = _RAND_3932[7:0];
  _RAND_3933 = {1{`RANDOM}};
  lineBuffer_3926 = _RAND_3933[7:0];
  _RAND_3934 = {1{`RANDOM}};
  lineBuffer_3927 = _RAND_3934[7:0];
  _RAND_3935 = {1{`RANDOM}};
  lineBuffer_3928 = _RAND_3935[7:0];
  _RAND_3936 = {1{`RANDOM}};
  lineBuffer_3929 = _RAND_3936[7:0];
  _RAND_3937 = {1{`RANDOM}};
  lineBuffer_3930 = _RAND_3937[7:0];
  _RAND_3938 = {1{`RANDOM}};
  lineBuffer_3931 = _RAND_3938[7:0];
  _RAND_3939 = {1{`RANDOM}};
  lineBuffer_3932 = _RAND_3939[7:0];
  _RAND_3940 = {1{`RANDOM}};
  lineBuffer_3933 = _RAND_3940[7:0];
  _RAND_3941 = {1{`RANDOM}};
  lineBuffer_3934 = _RAND_3941[7:0];
  _RAND_3942 = {1{`RANDOM}};
  lineBuffer_3935 = _RAND_3942[7:0];
  _RAND_3943 = {1{`RANDOM}};
  lineBuffer_3936 = _RAND_3943[7:0];
  _RAND_3944 = {1{`RANDOM}};
  lineBuffer_3937 = _RAND_3944[7:0];
  _RAND_3945 = {1{`RANDOM}};
  lineBuffer_3938 = _RAND_3945[7:0];
  _RAND_3946 = {1{`RANDOM}};
  lineBuffer_3939 = _RAND_3946[7:0];
  _RAND_3947 = {1{`RANDOM}};
  lineBuffer_3940 = _RAND_3947[7:0];
  _RAND_3948 = {1{`RANDOM}};
  lineBuffer_3941 = _RAND_3948[7:0];
  _RAND_3949 = {1{`RANDOM}};
  lineBuffer_3942 = _RAND_3949[7:0];
  _RAND_3950 = {1{`RANDOM}};
  lineBuffer_3943 = _RAND_3950[7:0];
  _RAND_3951 = {1{`RANDOM}};
  lineBuffer_3944 = _RAND_3951[7:0];
  _RAND_3952 = {1{`RANDOM}};
  lineBuffer_3945 = _RAND_3952[7:0];
  _RAND_3953 = {1{`RANDOM}};
  lineBuffer_3946 = _RAND_3953[7:0];
  _RAND_3954 = {1{`RANDOM}};
  lineBuffer_3947 = _RAND_3954[7:0];
  _RAND_3955 = {1{`RANDOM}};
  lineBuffer_3948 = _RAND_3955[7:0];
  _RAND_3956 = {1{`RANDOM}};
  lineBuffer_3949 = _RAND_3956[7:0];
  _RAND_3957 = {1{`RANDOM}};
  lineBuffer_3950 = _RAND_3957[7:0];
  _RAND_3958 = {1{`RANDOM}};
  lineBuffer_3951 = _RAND_3958[7:0];
  _RAND_3959 = {1{`RANDOM}};
  lineBuffer_3952 = _RAND_3959[7:0];
  _RAND_3960 = {1{`RANDOM}};
  lineBuffer_3953 = _RAND_3960[7:0];
  _RAND_3961 = {1{`RANDOM}};
  lineBuffer_3954 = _RAND_3961[7:0];
  _RAND_3962 = {1{`RANDOM}};
  lineBuffer_3955 = _RAND_3962[7:0];
  _RAND_3963 = {1{`RANDOM}};
  lineBuffer_3956 = _RAND_3963[7:0];
  _RAND_3964 = {1{`RANDOM}};
  lineBuffer_3957 = _RAND_3964[7:0];
  _RAND_3965 = {1{`RANDOM}};
  lineBuffer_3958 = _RAND_3965[7:0];
  _RAND_3966 = {1{`RANDOM}};
  lineBuffer_3959 = _RAND_3966[7:0];
  _RAND_3967 = {1{`RANDOM}};
  lineBuffer_3960 = _RAND_3967[7:0];
  _RAND_3968 = {1{`RANDOM}};
  lineBuffer_3961 = _RAND_3968[7:0];
  _RAND_3969 = {1{`RANDOM}};
  lineBuffer_3962 = _RAND_3969[7:0];
  _RAND_3970 = {1{`RANDOM}};
  lineBuffer_3963 = _RAND_3970[7:0];
  _RAND_3971 = {1{`RANDOM}};
  lineBuffer_3964 = _RAND_3971[7:0];
  _RAND_3972 = {1{`RANDOM}};
  lineBuffer_3965 = _RAND_3972[7:0];
  _RAND_3973 = {1{`RANDOM}};
  lineBuffer_3966 = _RAND_3973[7:0];
  _RAND_3974 = {1{`RANDOM}};
  lineBuffer_3967 = _RAND_3974[7:0];
  _RAND_3975 = {1{`RANDOM}};
  lineBuffer_3968 = _RAND_3975[7:0];
  _RAND_3976 = {1{`RANDOM}};
  lineBuffer_3969 = _RAND_3976[7:0];
  _RAND_3977 = {1{`RANDOM}};
  lineBuffer_3970 = _RAND_3977[7:0];
  _RAND_3978 = {1{`RANDOM}};
  lineBuffer_3971 = _RAND_3978[7:0];
  _RAND_3979 = {1{`RANDOM}};
  lineBuffer_3972 = _RAND_3979[7:0];
  _RAND_3980 = {1{`RANDOM}};
  lineBuffer_3973 = _RAND_3980[7:0];
  _RAND_3981 = {1{`RANDOM}};
  lineBuffer_3974 = _RAND_3981[7:0];
  _RAND_3982 = {1{`RANDOM}};
  lineBuffer_3975 = _RAND_3982[7:0];
  _RAND_3983 = {1{`RANDOM}};
  lineBuffer_3976 = _RAND_3983[7:0];
  _RAND_3984 = {1{`RANDOM}};
  lineBuffer_3977 = _RAND_3984[7:0];
  _RAND_3985 = {1{`RANDOM}};
  lineBuffer_3978 = _RAND_3985[7:0];
  _RAND_3986 = {1{`RANDOM}};
  lineBuffer_3979 = _RAND_3986[7:0];
  _RAND_3987 = {1{`RANDOM}};
  lineBuffer_3980 = _RAND_3987[7:0];
  _RAND_3988 = {1{`RANDOM}};
  lineBuffer_3981 = _RAND_3988[7:0];
  _RAND_3989 = {1{`RANDOM}};
  lineBuffer_3982 = _RAND_3989[7:0];
  _RAND_3990 = {1{`RANDOM}};
  lineBuffer_3983 = _RAND_3990[7:0];
  _RAND_3991 = {1{`RANDOM}};
  lineBuffer_3984 = _RAND_3991[7:0];
  _RAND_3992 = {1{`RANDOM}};
  lineBuffer_3985 = _RAND_3992[7:0];
  _RAND_3993 = {1{`RANDOM}};
  lineBuffer_3986 = _RAND_3993[7:0];
  _RAND_3994 = {1{`RANDOM}};
  lineBuffer_3987 = _RAND_3994[7:0];
  _RAND_3995 = {1{`RANDOM}};
  lineBuffer_3988 = _RAND_3995[7:0];
  _RAND_3996 = {1{`RANDOM}};
  lineBuffer_3989 = _RAND_3996[7:0];
  _RAND_3997 = {1{`RANDOM}};
  lineBuffer_3990 = _RAND_3997[7:0];
  _RAND_3998 = {1{`RANDOM}};
  lineBuffer_3991 = _RAND_3998[7:0];
  _RAND_3999 = {1{`RANDOM}};
  lineBuffer_3992 = _RAND_3999[7:0];
  _RAND_4000 = {1{`RANDOM}};
  lineBuffer_3993 = _RAND_4000[7:0];
  _RAND_4001 = {1{`RANDOM}};
  lineBuffer_3994 = _RAND_4001[7:0];
  _RAND_4002 = {1{`RANDOM}};
  lineBuffer_3995 = _RAND_4002[7:0];
  _RAND_4003 = {1{`RANDOM}};
  lineBuffer_3996 = _RAND_4003[7:0];
  _RAND_4004 = {1{`RANDOM}};
  lineBuffer_3997 = _RAND_4004[7:0];
  _RAND_4005 = {1{`RANDOM}};
  lineBuffer_3998 = _RAND_4005[7:0];
  _RAND_4006 = {1{`RANDOM}};
  lineBuffer_3999 = _RAND_4006[7:0];
  _RAND_4007 = {1{`RANDOM}};
  lineBuffer_4000 = _RAND_4007[7:0];
  _RAND_4008 = {1{`RANDOM}};
  lineBuffer_4001 = _RAND_4008[7:0];
  _RAND_4009 = {1{`RANDOM}};
  lineBuffer_4002 = _RAND_4009[7:0];
  _RAND_4010 = {1{`RANDOM}};
  lineBuffer_4003 = _RAND_4010[7:0];
  _RAND_4011 = {1{`RANDOM}};
  lineBuffer_4004 = _RAND_4011[7:0];
  _RAND_4012 = {1{`RANDOM}};
  lineBuffer_4005 = _RAND_4012[7:0];
  _RAND_4013 = {1{`RANDOM}};
  lineBuffer_4006 = _RAND_4013[7:0];
  _RAND_4014 = {1{`RANDOM}};
  lineBuffer_4007 = _RAND_4014[7:0];
  _RAND_4015 = {1{`RANDOM}};
  lineBuffer_4008 = _RAND_4015[7:0];
  _RAND_4016 = {1{`RANDOM}};
  lineBuffer_4009 = _RAND_4016[7:0];
  _RAND_4017 = {1{`RANDOM}};
  lineBuffer_4010 = _RAND_4017[7:0];
  _RAND_4018 = {1{`RANDOM}};
  lineBuffer_4011 = _RAND_4018[7:0];
  _RAND_4019 = {1{`RANDOM}};
  lineBuffer_4012 = _RAND_4019[7:0];
  _RAND_4020 = {1{`RANDOM}};
  lineBuffer_4013 = _RAND_4020[7:0];
  _RAND_4021 = {1{`RANDOM}};
  lineBuffer_4014 = _RAND_4021[7:0];
  _RAND_4022 = {1{`RANDOM}};
  lineBuffer_4015 = _RAND_4022[7:0];
  _RAND_4023 = {1{`RANDOM}};
  lineBuffer_4016 = _RAND_4023[7:0];
  _RAND_4024 = {1{`RANDOM}};
  lineBuffer_4017 = _RAND_4024[7:0];
  _RAND_4025 = {1{`RANDOM}};
  lineBuffer_4018 = _RAND_4025[7:0];
  _RAND_4026 = {1{`RANDOM}};
  lineBuffer_4019 = _RAND_4026[7:0];
  _RAND_4027 = {1{`RANDOM}};
  lineBuffer_4020 = _RAND_4027[7:0];
  _RAND_4028 = {1{`RANDOM}};
  lineBuffer_4021 = _RAND_4028[7:0];
  _RAND_4029 = {1{`RANDOM}};
  lineBuffer_4022 = _RAND_4029[7:0];
  _RAND_4030 = {1{`RANDOM}};
  lineBuffer_4023 = _RAND_4030[7:0];
  _RAND_4031 = {1{`RANDOM}};
  lineBuffer_4024 = _RAND_4031[7:0];
  _RAND_4032 = {1{`RANDOM}};
  lineBuffer_4025 = _RAND_4032[7:0];
  _RAND_4033 = {1{`RANDOM}};
  lineBuffer_4026 = _RAND_4033[7:0];
  _RAND_4034 = {1{`RANDOM}};
  lineBuffer_4027 = _RAND_4034[7:0];
  _RAND_4035 = {1{`RANDOM}};
  lineBuffer_4028 = _RAND_4035[7:0];
  _RAND_4036 = {1{`RANDOM}};
  lineBuffer_4029 = _RAND_4036[7:0];
  _RAND_4037 = {1{`RANDOM}};
  lineBuffer_4030 = _RAND_4037[7:0];
  _RAND_4038 = {1{`RANDOM}};
  lineBuffer_4031 = _RAND_4038[7:0];
  _RAND_4039 = {1{`RANDOM}};
  lineBuffer_4032 = _RAND_4039[7:0];
  _RAND_4040 = {1{`RANDOM}};
  lineBuffer_4033 = _RAND_4040[7:0];
  _RAND_4041 = {1{`RANDOM}};
  lineBuffer_4034 = _RAND_4041[7:0];
  _RAND_4042 = {1{`RANDOM}};
  lineBuffer_4035 = _RAND_4042[7:0];
  _RAND_4043 = {1{`RANDOM}};
  lineBuffer_4036 = _RAND_4043[7:0];
  _RAND_4044 = {1{`RANDOM}};
  lineBuffer_4037 = _RAND_4044[7:0];
  _RAND_4045 = {1{`RANDOM}};
  lineBuffer_4038 = _RAND_4045[7:0];
  _RAND_4046 = {1{`RANDOM}};
  lineBuffer_4039 = _RAND_4046[7:0];
  _RAND_4047 = {1{`RANDOM}};
  lineBuffer_4040 = _RAND_4047[7:0];
  _RAND_4048 = {1{`RANDOM}};
  lineBuffer_4041 = _RAND_4048[7:0];
  _RAND_4049 = {1{`RANDOM}};
  lineBuffer_4042 = _RAND_4049[7:0];
  _RAND_4050 = {1{`RANDOM}};
  lineBuffer_4043 = _RAND_4050[7:0];
  _RAND_4051 = {1{`RANDOM}};
  lineBuffer_4044 = _RAND_4051[7:0];
  _RAND_4052 = {1{`RANDOM}};
  lineBuffer_4045 = _RAND_4052[7:0];
  _RAND_4053 = {1{`RANDOM}};
  lineBuffer_4046 = _RAND_4053[7:0];
  _RAND_4054 = {1{`RANDOM}};
  lineBuffer_4047 = _RAND_4054[7:0];
  _RAND_4055 = {1{`RANDOM}};
  lineBuffer_4048 = _RAND_4055[7:0];
  _RAND_4056 = {1{`RANDOM}};
  lineBuffer_4049 = _RAND_4056[7:0];
  _RAND_4057 = {1{`RANDOM}};
  lineBuffer_4050 = _RAND_4057[7:0];
  _RAND_4058 = {1{`RANDOM}};
  lineBuffer_4051 = _RAND_4058[7:0];
  _RAND_4059 = {1{`RANDOM}};
  lineBuffer_4052 = _RAND_4059[7:0];
  _RAND_4060 = {1{`RANDOM}};
  lineBuffer_4053 = _RAND_4060[7:0];
  _RAND_4061 = {1{`RANDOM}};
  lineBuffer_4054 = _RAND_4061[7:0];
  _RAND_4062 = {1{`RANDOM}};
  lineBuffer_4055 = _RAND_4062[7:0];
  _RAND_4063 = {1{`RANDOM}};
  lineBuffer_4056 = _RAND_4063[7:0];
  _RAND_4064 = {1{`RANDOM}};
  lineBuffer_4057 = _RAND_4064[7:0];
  _RAND_4065 = {1{`RANDOM}};
  lineBuffer_4058 = _RAND_4065[7:0];
  _RAND_4066 = {1{`RANDOM}};
  lineBuffer_4059 = _RAND_4066[7:0];
  _RAND_4067 = {1{`RANDOM}};
  lineBuffer_4060 = _RAND_4067[7:0];
  _RAND_4068 = {1{`RANDOM}};
  lineBuffer_4061 = _RAND_4068[7:0];
  _RAND_4069 = {1{`RANDOM}};
  lineBuffer_4062 = _RAND_4069[7:0];
  _RAND_4070 = {1{`RANDOM}};
  lineBuffer_4063 = _RAND_4070[7:0];
  _RAND_4071 = {1{`RANDOM}};
  lineBuffer_4064 = _RAND_4071[7:0];
  _RAND_4072 = {1{`RANDOM}};
  lineBuffer_4065 = _RAND_4072[7:0];
  _RAND_4073 = {1{`RANDOM}};
  lineBuffer_4066 = _RAND_4073[7:0];
  _RAND_4074 = {1{`RANDOM}};
  lineBuffer_4067 = _RAND_4074[7:0];
  _RAND_4075 = {1{`RANDOM}};
  lineBuffer_4068 = _RAND_4075[7:0];
  _RAND_4076 = {1{`RANDOM}};
  lineBuffer_4069 = _RAND_4076[7:0];
  _RAND_4077 = {1{`RANDOM}};
  lineBuffer_4070 = _RAND_4077[7:0];
  _RAND_4078 = {1{`RANDOM}};
  lineBuffer_4071 = _RAND_4078[7:0];
  _RAND_4079 = {1{`RANDOM}};
  lineBuffer_4072 = _RAND_4079[7:0];
  _RAND_4080 = {1{`RANDOM}};
  lineBuffer_4073 = _RAND_4080[7:0];
  _RAND_4081 = {1{`RANDOM}};
  lineBuffer_4074 = _RAND_4081[7:0];
  _RAND_4082 = {1{`RANDOM}};
  lineBuffer_4075 = _RAND_4082[7:0];
  _RAND_4083 = {1{`RANDOM}};
  lineBuffer_4076 = _RAND_4083[7:0];
  _RAND_4084 = {1{`RANDOM}};
  lineBuffer_4077 = _RAND_4084[7:0];
  _RAND_4085 = {1{`RANDOM}};
  lineBuffer_4078 = _RAND_4085[7:0];
  _RAND_4086 = {1{`RANDOM}};
  lineBuffer_4079 = _RAND_4086[7:0];
  _RAND_4087 = {1{`RANDOM}};
  lineBuffer_4080 = _RAND_4087[7:0];
  _RAND_4088 = {1{`RANDOM}};
  lineBuffer_4081 = _RAND_4088[7:0];
  _RAND_4089 = {1{`RANDOM}};
  lineBuffer_4082 = _RAND_4089[7:0];
  _RAND_4090 = {1{`RANDOM}};
  lineBuffer_4083 = _RAND_4090[7:0];
  _RAND_4091 = {1{`RANDOM}};
  lineBuffer_4084 = _RAND_4091[7:0];
  _RAND_4092 = {1{`RANDOM}};
  lineBuffer_4085 = _RAND_4092[7:0];
  _RAND_4093 = {1{`RANDOM}};
  lineBuffer_4086 = _RAND_4093[7:0];
  _RAND_4094 = {1{`RANDOM}};
  lineBuffer_4087 = _RAND_4094[7:0];
  _RAND_4095 = {1{`RANDOM}};
  lineBuffer_4088 = _RAND_4095[7:0];
  _RAND_4096 = {1{`RANDOM}};
  lineBuffer_4089 = _RAND_4096[7:0];
  _RAND_4097 = {1{`RANDOM}};
  lineBuffer_4090 = _RAND_4097[7:0];
  _RAND_4098 = {1{`RANDOM}};
  lineBuffer_4091 = _RAND_4098[7:0];
  _RAND_4099 = {1{`RANDOM}};
  lineBuffer_4092 = _RAND_4099[7:0];
  _RAND_4100 = {1{`RANDOM}};
  lineBuffer_4093 = _RAND_4100[7:0];
  _RAND_4101 = {1{`RANDOM}};
  lineBuffer_4094 = _RAND_4101[7:0];
  _RAND_4102 = {1{`RANDOM}};
  lineBuffer_4095 = _RAND_4102[7:0];
  _RAND_4103 = {1{`RANDOM}};
  lineBuffer_4096 = _RAND_4103[7:0];
  _RAND_4104 = {1{`RANDOM}};
  lineBuffer_4097 = _RAND_4104[7:0];
  _RAND_4105 = {1{`RANDOM}};
  lineBuffer_4098 = _RAND_4105[7:0];
  _RAND_4106 = {1{`RANDOM}};
  lineBuffer_4099 = _RAND_4106[7:0];
  _RAND_4107 = {1{`RANDOM}};
  lineBuffer_4100 = _RAND_4107[7:0];
  _RAND_4108 = {1{`RANDOM}};
  lineBuffer_4101 = _RAND_4108[7:0];
  _RAND_4109 = {1{`RANDOM}};
  lineBuffer_4102 = _RAND_4109[7:0];
  _RAND_4110 = {1{`RANDOM}};
  lineBuffer_4103 = _RAND_4110[7:0];
  _RAND_4111 = {1{`RANDOM}};
  lineBuffer_4104 = _RAND_4111[7:0];
  _RAND_4112 = {1{`RANDOM}};
  lineBuffer_4105 = _RAND_4112[7:0];
  _RAND_4113 = {1{`RANDOM}};
  lineBuffer_4106 = _RAND_4113[7:0];
  _RAND_4114 = {1{`RANDOM}};
  lineBuffer_4107 = _RAND_4114[7:0];
  _RAND_4115 = {1{`RANDOM}};
  lineBuffer_4108 = _RAND_4115[7:0];
  _RAND_4116 = {1{`RANDOM}};
  lineBuffer_4109 = _RAND_4116[7:0];
  _RAND_4117 = {1{`RANDOM}};
  lineBuffer_4110 = _RAND_4117[7:0];
  _RAND_4118 = {1{`RANDOM}};
  lineBuffer_4111 = _RAND_4118[7:0];
  _RAND_4119 = {1{`RANDOM}};
  lineBuffer_4112 = _RAND_4119[7:0];
  _RAND_4120 = {1{`RANDOM}};
  lineBuffer_4113 = _RAND_4120[7:0];
  _RAND_4121 = {1{`RANDOM}};
  lineBuffer_4114 = _RAND_4121[7:0];
  _RAND_4122 = {1{`RANDOM}};
  lineBuffer_4115 = _RAND_4122[7:0];
  _RAND_4123 = {1{`RANDOM}};
  lineBuffer_4116 = _RAND_4123[7:0];
  _RAND_4124 = {1{`RANDOM}};
  lineBuffer_4117 = _RAND_4124[7:0];
  _RAND_4125 = {1{`RANDOM}};
  lineBuffer_4118 = _RAND_4125[7:0];
  _RAND_4126 = {1{`RANDOM}};
  lineBuffer_4119 = _RAND_4126[7:0];
  _RAND_4127 = {1{`RANDOM}};
  lineBuffer_4120 = _RAND_4127[7:0];
  _RAND_4128 = {1{`RANDOM}};
  lineBuffer_4121 = _RAND_4128[7:0];
  _RAND_4129 = {1{`RANDOM}};
  lineBuffer_4122 = _RAND_4129[7:0];
  _RAND_4130 = {1{`RANDOM}};
  lineBuffer_4123 = _RAND_4130[7:0];
  _RAND_4131 = {1{`RANDOM}};
  lineBuffer_4124 = _RAND_4131[7:0];
  _RAND_4132 = {1{`RANDOM}};
  lineBuffer_4125 = _RAND_4132[7:0];
  _RAND_4133 = {1{`RANDOM}};
  lineBuffer_4126 = _RAND_4133[7:0];
  _RAND_4134 = {1{`RANDOM}};
  lineBuffer_4127 = _RAND_4134[7:0];
  _RAND_4135 = {1{`RANDOM}};
  lineBuffer_4128 = _RAND_4135[7:0];
  _RAND_4136 = {1{`RANDOM}};
  lineBuffer_4129 = _RAND_4136[7:0];
  _RAND_4137 = {1{`RANDOM}};
  lineBuffer_4130 = _RAND_4137[7:0];
  _RAND_4138 = {1{`RANDOM}};
  lineBuffer_4131 = _RAND_4138[7:0];
  _RAND_4139 = {1{`RANDOM}};
  lineBuffer_4132 = _RAND_4139[7:0];
  _RAND_4140 = {1{`RANDOM}};
  lineBuffer_4133 = _RAND_4140[7:0];
  _RAND_4141 = {1{`RANDOM}};
  lineBuffer_4134 = _RAND_4141[7:0];
  _RAND_4142 = {1{`RANDOM}};
  lineBuffer_4135 = _RAND_4142[7:0];
  _RAND_4143 = {1{`RANDOM}};
  lineBuffer_4136 = _RAND_4143[7:0];
  _RAND_4144 = {1{`RANDOM}};
  lineBuffer_4137 = _RAND_4144[7:0];
  _RAND_4145 = {1{`RANDOM}};
  lineBuffer_4138 = _RAND_4145[7:0];
  _RAND_4146 = {1{`RANDOM}};
  lineBuffer_4139 = _RAND_4146[7:0];
  _RAND_4147 = {1{`RANDOM}};
  lineBuffer_4140 = _RAND_4147[7:0];
  _RAND_4148 = {1{`RANDOM}};
  lineBuffer_4141 = _RAND_4148[7:0];
  _RAND_4149 = {1{`RANDOM}};
  lineBuffer_4142 = _RAND_4149[7:0];
  _RAND_4150 = {1{`RANDOM}};
  lineBuffer_4143 = _RAND_4150[7:0];
  _RAND_4151 = {1{`RANDOM}};
  lineBuffer_4144 = _RAND_4151[7:0];
  _RAND_4152 = {1{`RANDOM}};
  lineBuffer_4145 = _RAND_4152[7:0];
  _RAND_4153 = {1{`RANDOM}};
  lineBuffer_4146 = _RAND_4153[7:0];
  _RAND_4154 = {1{`RANDOM}};
  lineBuffer_4147 = _RAND_4154[7:0];
  _RAND_4155 = {1{`RANDOM}};
  lineBuffer_4148 = _RAND_4155[7:0];
  _RAND_4156 = {1{`RANDOM}};
  lineBuffer_4149 = _RAND_4156[7:0];
  _RAND_4157 = {1{`RANDOM}};
  lineBuffer_4150 = _RAND_4157[7:0];
  _RAND_4158 = {1{`RANDOM}};
  lineBuffer_4151 = _RAND_4158[7:0];
  _RAND_4159 = {1{`RANDOM}};
  lineBuffer_4152 = _RAND_4159[7:0];
  _RAND_4160 = {1{`RANDOM}};
  lineBuffer_4153 = _RAND_4160[7:0];
  _RAND_4161 = {1{`RANDOM}};
  lineBuffer_4154 = _RAND_4161[7:0];
  _RAND_4162 = {1{`RANDOM}};
  lineBuffer_4155 = _RAND_4162[7:0];
  _RAND_4163 = {1{`RANDOM}};
  lineBuffer_4156 = _RAND_4163[7:0];
  _RAND_4164 = {1{`RANDOM}};
  lineBuffer_4157 = _RAND_4164[7:0];
  _RAND_4165 = {1{`RANDOM}};
  lineBuffer_4158 = _RAND_4165[7:0];
  _RAND_4166 = {1{`RANDOM}};
  lineBuffer_4159 = _RAND_4166[7:0];
  _RAND_4167 = {1{`RANDOM}};
  lineBuffer_4160 = _RAND_4167[7:0];
  _RAND_4168 = {1{`RANDOM}};
  lineBuffer_4161 = _RAND_4168[7:0];
  _RAND_4169 = {1{`RANDOM}};
  lineBuffer_4162 = _RAND_4169[7:0];
  _RAND_4170 = {1{`RANDOM}};
  lineBuffer_4163 = _RAND_4170[7:0];
  _RAND_4171 = {1{`RANDOM}};
  lineBuffer_4164 = _RAND_4171[7:0];
  _RAND_4172 = {1{`RANDOM}};
  lineBuffer_4165 = _RAND_4172[7:0];
  _RAND_4173 = {1{`RANDOM}};
  lineBuffer_4166 = _RAND_4173[7:0];
  _RAND_4174 = {1{`RANDOM}};
  lineBuffer_4167 = _RAND_4174[7:0];
  _RAND_4175 = {1{`RANDOM}};
  lineBuffer_4168 = _RAND_4175[7:0];
  _RAND_4176 = {1{`RANDOM}};
  lineBuffer_4169 = _RAND_4176[7:0];
  _RAND_4177 = {1{`RANDOM}};
  lineBuffer_4170 = _RAND_4177[7:0];
  _RAND_4178 = {1{`RANDOM}};
  lineBuffer_4171 = _RAND_4178[7:0];
  _RAND_4179 = {1{`RANDOM}};
  lineBuffer_4172 = _RAND_4179[7:0];
  _RAND_4180 = {1{`RANDOM}};
  lineBuffer_4173 = _RAND_4180[7:0];
  _RAND_4181 = {1{`RANDOM}};
  lineBuffer_4174 = _RAND_4181[7:0];
  _RAND_4182 = {1{`RANDOM}};
  lineBuffer_4175 = _RAND_4182[7:0];
  _RAND_4183 = {1{`RANDOM}};
  lineBuffer_4176 = _RAND_4183[7:0];
  _RAND_4184 = {1{`RANDOM}};
  lineBuffer_4177 = _RAND_4184[7:0];
  _RAND_4185 = {1{`RANDOM}};
  lineBuffer_4178 = _RAND_4185[7:0];
  _RAND_4186 = {1{`RANDOM}};
  lineBuffer_4179 = _RAND_4186[7:0];
  _RAND_4187 = {1{`RANDOM}};
  lineBuffer_4180 = _RAND_4187[7:0];
  _RAND_4188 = {1{`RANDOM}};
  lineBuffer_4181 = _RAND_4188[7:0];
  _RAND_4189 = {1{`RANDOM}};
  lineBuffer_4182 = _RAND_4189[7:0];
  _RAND_4190 = {1{`RANDOM}};
  lineBuffer_4183 = _RAND_4190[7:0];
  _RAND_4191 = {1{`RANDOM}};
  lineBuffer_4184 = _RAND_4191[7:0];
  _RAND_4192 = {1{`RANDOM}};
  lineBuffer_4185 = _RAND_4192[7:0];
  _RAND_4193 = {1{`RANDOM}};
  lineBuffer_4186 = _RAND_4193[7:0];
  _RAND_4194 = {1{`RANDOM}};
  lineBuffer_4187 = _RAND_4194[7:0];
  _RAND_4195 = {1{`RANDOM}};
  lineBuffer_4188 = _RAND_4195[7:0];
  _RAND_4196 = {1{`RANDOM}};
  lineBuffer_4189 = _RAND_4196[7:0];
  _RAND_4197 = {1{`RANDOM}};
  lineBuffer_4190 = _RAND_4197[7:0];
  _RAND_4198 = {1{`RANDOM}};
  lineBuffer_4191 = _RAND_4198[7:0];
  _RAND_4199 = {1{`RANDOM}};
  lineBuffer_4192 = _RAND_4199[7:0];
  _RAND_4200 = {1{`RANDOM}};
  lineBuffer_4193 = _RAND_4200[7:0];
  _RAND_4201 = {1{`RANDOM}};
  lineBuffer_4194 = _RAND_4201[7:0];
  _RAND_4202 = {1{`RANDOM}};
  lineBuffer_4195 = _RAND_4202[7:0];
  _RAND_4203 = {1{`RANDOM}};
  lineBuffer_4196 = _RAND_4203[7:0];
  _RAND_4204 = {1{`RANDOM}};
  lineBuffer_4197 = _RAND_4204[7:0];
  _RAND_4205 = {1{`RANDOM}};
  lineBuffer_4198 = _RAND_4205[7:0];
  _RAND_4206 = {1{`RANDOM}};
  lineBuffer_4199 = _RAND_4206[7:0];
  _RAND_4207 = {1{`RANDOM}};
  lineBuffer_4200 = _RAND_4207[7:0];
  _RAND_4208 = {1{`RANDOM}};
  lineBuffer_4201 = _RAND_4208[7:0];
  _RAND_4209 = {1{`RANDOM}};
  lineBuffer_4202 = _RAND_4209[7:0];
  _RAND_4210 = {1{`RANDOM}};
  lineBuffer_4203 = _RAND_4210[7:0];
  _RAND_4211 = {1{`RANDOM}};
  lineBuffer_4204 = _RAND_4211[7:0];
  _RAND_4212 = {1{`RANDOM}};
  lineBuffer_4205 = _RAND_4212[7:0];
  _RAND_4213 = {1{`RANDOM}};
  lineBuffer_4206 = _RAND_4213[7:0];
  _RAND_4214 = {1{`RANDOM}};
  lineBuffer_4207 = _RAND_4214[7:0];
  _RAND_4215 = {1{`RANDOM}};
  lineBuffer_4208 = _RAND_4215[7:0];
  _RAND_4216 = {1{`RANDOM}};
  lineBuffer_4209 = _RAND_4216[7:0];
  _RAND_4217 = {1{`RANDOM}};
  lineBuffer_4210 = _RAND_4217[7:0];
  _RAND_4218 = {1{`RANDOM}};
  lineBuffer_4211 = _RAND_4218[7:0];
  _RAND_4219 = {1{`RANDOM}};
  lineBuffer_4212 = _RAND_4219[7:0];
  _RAND_4220 = {1{`RANDOM}};
  lineBuffer_4213 = _RAND_4220[7:0];
  _RAND_4221 = {1{`RANDOM}};
  lineBuffer_4214 = _RAND_4221[7:0];
  _RAND_4222 = {1{`RANDOM}};
  lineBuffer_4215 = _RAND_4222[7:0];
  _RAND_4223 = {1{`RANDOM}};
  lineBuffer_4216 = _RAND_4223[7:0];
  _RAND_4224 = {1{`RANDOM}};
  lineBuffer_4217 = _RAND_4224[7:0];
  _RAND_4225 = {1{`RANDOM}};
  lineBuffer_4218 = _RAND_4225[7:0];
  _RAND_4226 = {1{`RANDOM}};
  lineBuffer_4219 = _RAND_4226[7:0];
  _RAND_4227 = {1{`RANDOM}};
  lineBuffer_4220 = _RAND_4227[7:0];
  _RAND_4228 = {1{`RANDOM}};
  lineBuffer_4221 = _RAND_4228[7:0];
  _RAND_4229 = {1{`RANDOM}};
  lineBuffer_4222 = _RAND_4229[7:0];
  _RAND_4230 = {1{`RANDOM}};
  lineBuffer_4223 = _RAND_4230[7:0];
  _RAND_4231 = {1{`RANDOM}};
  lineBuffer_4224 = _RAND_4231[7:0];
  _RAND_4232 = {1{`RANDOM}};
  lineBuffer_4225 = _RAND_4232[7:0];
  _RAND_4233 = {1{`RANDOM}};
  lineBuffer_4226 = _RAND_4233[7:0];
  _RAND_4234 = {1{`RANDOM}};
  lineBuffer_4227 = _RAND_4234[7:0];
  _RAND_4235 = {1{`RANDOM}};
  lineBuffer_4228 = _RAND_4235[7:0];
  _RAND_4236 = {1{`RANDOM}};
  lineBuffer_4229 = _RAND_4236[7:0];
  _RAND_4237 = {1{`RANDOM}};
  lineBuffer_4230 = _RAND_4237[7:0];
  _RAND_4238 = {1{`RANDOM}};
  lineBuffer_4231 = _RAND_4238[7:0];
  _RAND_4239 = {1{`RANDOM}};
  lineBuffer_4232 = _RAND_4239[7:0];
  _RAND_4240 = {1{`RANDOM}};
  lineBuffer_4233 = _RAND_4240[7:0];
  _RAND_4241 = {1{`RANDOM}};
  lineBuffer_4234 = _RAND_4241[7:0];
  _RAND_4242 = {1{`RANDOM}};
  lineBuffer_4235 = _RAND_4242[7:0];
  _RAND_4243 = {1{`RANDOM}};
  lineBuffer_4236 = _RAND_4243[7:0];
  _RAND_4244 = {1{`RANDOM}};
  lineBuffer_4237 = _RAND_4244[7:0];
  _RAND_4245 = {1{`RANDOM}};
  lineBuffer_4238 = _RAND_4245[7:0];
  _RAND_4246 = {1{`RANDOM}};
  lineBuffer_4239 = _RAND_4246[7:0];
  _RAND_4247 = {1{`RANDOM}};
  lineBuffer_4240 = _RAND_4247[7:0];
  _RAND_4248 = {1{`RANDOM}};
  lineBuffer_4241 = _RAND_4248[7:0];
  _RAND_4249 = {1{`RANDOM}};
  lineBuffer_4242 = _RAND_4249[7:0];
  _RAND_4250 = {1{`RANDOM}};
  lineBuffer_4243 = _RAND_4250[7:0];
  _RAND_4251 = {1{`RANDOM}};
  lineBuffer_4244 = _RAND_4251[7:0];
  _RAND_4252 = {1{`RANDOM}};
  lineBuffer_4245 = _RAND_4252[7:0];
  _RAND_4253 = {1{`RANDOM}};
  lineBuffer_4246 = _RAND_4253[7:0];
  _RAND_4254 = {1{`RANDOM}};
  lineBuffer_4247 = _RAND_4254[7:0];
  _RAND_4255 = {1{`RANDOM}};
  lineBuffer_4248 = _RAND_4255[7:0];
  _RAND_4256 = {1{`RANDOM}};
  lineBuffer_4249 = _RAND_4256[7:0];
  _RAND_4257 = {1{`RANDOM}};
  lineBuffer_4250 = _RAND_4257[7:0];
  _RAND_4258 = {1{`RANDOM}};
  lineBuffer_4251 = _RAND_4258[7:0];
  _RAND_4259 = {1{`RANDOM}};
  lineBuffer_4252 = _RAND_4259[7:0];
  _RAND_4260 = {1{`RANDOM}};
  lineBuffer_4253 = _RAND_4260[7:0];
  _RAND_4261 = {1{`RANDOM}};
  lineBuffer_4254 = _RAND_4261[7:0];
  _RAND_4262 = {1{`RANDOM}};
  lineBuffer_4255 = _RAND_4262[7:0];
  _RAND_4263 = {1{`RANDOM}};
  lineBuffer_4256 = _RAND_4263[7:0];
  _RAND_4264 = {1{`RANDOM}};
  lineBuffer_4257 = _RAND_4264[7:0];
  _RAND_4265 = {1{`RANDOM}};
  lineBuffer_4258 = _RAND_4265[7:0];
  _RAND_4266 = {1{`RANDOM}};
  lineBuffer_4259 = _RAND_4266[7:0];
  _RAND_4267 = {1{`RANDOM}};
  lineBuffer_4260 = _RAND_4267[7:0];
  _RAND_4268 = {1{`RANDOM}};
  lineBuffer_4261 = _RAND_4268[7:0];
  _RAND_4269 = {1{`RANDOM}};
  lineBuffer_4262 = _RAND_4269[7:0];
  _RAND_4270 = {1{`RANDOM}};
  lineBuffer_4263 = _RAND_4270[7:0];
  _RAND_4271 = {1{`RANDOM}};
  lineBuffer_4264 = _RAND_4271[7:0];
  _RAND_4272 = {1{`RANDOM}};
  lineBuffer_4265 = _RAND_4272[7:0];
  _RAND_4273 = {1{`RANDOM}};
  lineBuffer_4266 = _RAND_4273[7:0];
  _RAND_4274 = {1{`RANDOM}};
  lineBuffer_4267 = _RAND_4274[7:0];
  _RAND_4275 = {1{`RANDOM}};
  lineBuffer_4268 = _RAND_4275[7:0];
  _RAND_4276 = {1{`RANDOM}};
  lineBuffer_4269 = _RAND_4276[7:0];
  _RAND_4277 = {1{`RANDOM}};
  lineBuffer_4270 = _RAND_4277[7:0];
  _RAND_4278 = {1{`RANDOM}};
  lineBuffer_4271 = _RAND_4278[7:0];
  _RAND_4279 = {1{`RANDOM}};
  lineBuffer_4272 = _RAND_4279[7:0];
  _RAND_4280 = {1{`RANDOM}};
  lineBuffer_4273 = _RAND_4280[7:0];
  _RAND_4281 = {1{`RANDOM}};
  lineBuffer_4274 = _RAND_4281[7:0];
  _RAND_4282 = {1{`RANDOM}};
  lineBuffer_4275 = _RAND_4282[7:0];
  _RAND_4283 = {1{`RANDOM}};
  lineBuffer_4276 = _RAND_4283[7:0];
  _RAND_4284 = {1{`RANDOM}};
  lineBuffer_4277 = _RAND_4284[7:0];
  _RAND_4285 = {1{`RANDOM}};
  lineBuffer_4278 = _RAND_4285[7:0];
  _RAND_4286 = {1{`RANDOM}};
  lineBuffer_4279 = _RAND_4286[7:0];
  _RAND_4287 = {1{`RANDOM}};
  lineBuffer_4280 = _RAND_4287[7:0];
  _RAND_4288 = {1{`RANDOM}};
  lineBuffer_4281 = _RAND_4288[7:0];
  _RAND_4289 = {1{`RANDOM}};
  lineBuffer_4282 = _RAND_4289[7:0];
  _RAND_4290 = {1{`RANDOM}};
  lineBuffer_4283 = _RAND_4290[7:0];
  _RAND_4291 = {1{`RANDOM}};
  lineBuffer_4284 = _RAND_4291[7:0];
  _RAND_4292 = {1{`RANDOM}};
  lineBuffer_4285 = _RAND_4292[7:0];
  _RAND_4293 = {1{`RANDOM}};
  lineBuffer_4286 = _RAND_4293[7:0];
  _RAND_4294 = {1{`RANDOM}};
  lineBuffer_4287 = _RAND_4294[7:0];
  _RAND_4295 = {1{`RANDOM}};
  lineBuffer_4288 = _RAND_4295[7:0];
  _RAND_4296 = {1{`RANDOM}};
  lineBuffer_4289 = _RAND_4296[7:0];
  _RAND_4297 = {1{`RANDOM}};
  lineBuffer_4290 = _RAND_4297[7:0];
  _RAND_4298 = {1{`RANDOM}};
  lineBuffer_4291 = _RAND_4298[7:0];
  _RAND_4299 = {1{`RANDOM}};
  lineBuffer_4292 = _RAND_4299[7:0];
  _RAND_4300 = {1{`RANDOM}};
  lineBuffer_4293 = _RAND_4300[7:0];
  _RAND_4301 = {1{`RANDOM}};
  lineBuffer_4294 = _RAND_4301[7:0];
  _RAND_4302 = {1{`RANDOM}};
  lineBuffer_4295 = _RAND_4302[7:0];
  _RAND_4303 = {1{`RANDOM}};
  lineBuffer_4296 = _RAND_4303[7:0];
  _RAND_4304 = {1{`RANDOM}};
  lineBuffer_4297 = _RAND_4304[7:0];
  _RAND_4305 = {1{`RANDOM}};
  lineBuffer_4298 = _RAND_4305[7:0];
  _RAND_4306 = {1{`RANDOM}};
  lineBuffer_4299 = _RAND_4306[7:0];
  _RAND_4307 = {1{`RANDOM}};
  lineBuffer_4300 = _RAND_4307[7:0];
  _RAND_4308 = {1{`RANDOM}};
  lineBuffer_4301 = _RAND_4308[7:0];
  _RAND_4309 = {1{`RANDOM}};
  lineBuffer_4302 = _RAND_4309[7:0];
  _RAND_4310 = {1{`RANDOM}};
  lineBuffer_4303 = _RAND_4310[7:0];
  _RAND_4311 = {1{`RANDOM}};
  lineBuffer_4304 = _RAND_4311[7:0];
  _RAND_4312 = {1{`RANDOM}};
  lineBuffer_4305 = _RAND_4312[7:0];
  _RAND_4313 = {1{`RANDOM}};
  lineBuffer_4306 = _RAND_4313[7:0];
  _RAND_4314 = {1{`RANDOM}};
  lineBuffer_4307 = _RAND_4314[7:0];
  _RAND_4315 = {1{`RANDOM}};
  lineBuffer_4308 = _RAND_4315[7:0];
  _RAND_4316 = {1{`RANDOM}};
  lineBuffer_4309 = _RAND_4316[7:0];
  _RAND_4317 = {1{`RANDOM}};
  lineBuffer_4310 = _RAND_4317[7:0];
  _RAND_4318 = {1{`RANDOM}};
  lineBuffer_4311 = _RAND_4318[7:0];
  _RAND_4319 = {1{`RANDOM}};
  lineBuffer_4312 = _RAND_4319[7:0];
  _RAND_4320 = {1{`RANDOM}};
  lineBuffer_4313 = _RAND_4320[7:0];
  _RAND_4321 = {1{`RANDOM}};
  lineBuffer_4314 = _RAND_4321[7:0];
  _RAND_4322 = {1{`RANDOM}};
  lineBuffer_4315 = _RAND_4322[7:0];
  _RAND_4323 = {1{`RANDOM}};
  lineBuffer_4316 = _RAND_4323[7:0];
  _RAND_4324 = {1{`RANDOM}};
  lineBuffer_4317 = _RAND_4324[7:0];
  _RAND_4325 = {1{`RANDOM}};
  lineBuffer_4318 = _RAND_4325[7:0];
  _RAND_4326 = {1{`RANDOM}};
  lineBuffer_4319 = _RAND_4326[7:0];
  _RAND_4327 = {1{`RANDOM}};
  lineBuffer_4320 = _RAND_4327[7:0];
  _RAND_4328 = {1{`RANDOM}};
  lineBuffer_4321 = _RAND_4328[7:0];
  _RAND_4329 = {1{`RANDOM}};
  lineBuffer_4322 = _RAND_4329[7:0];
  _RAND_4330 = {1{`RANDOM}};
  lineBuffer_4323 = _RAND_4330[7:0];
  _RAND_4331 = {1{`RANDOM}};
  lineBuffer_4324 = _RAND_4331[7:0];
  _RAND_4332 = {1{`RANDOM}};
  lineBuffer_4325 = _RAND_4332[7:0];
  _RAND_4333 = {1{`RANDOM}};
  lineBuffer_4326 = _RAND_4333[7:0];
  _RAND_4334 = {1{`RANDOM}};
  lineBuffer_4327 = _RAND_4334[7:0];
  _RAND_4335 = {1{`RANDOM}};
  lineBuffer_4328 = _RAND_4335[7:0];
  _RAND_4336 = {1{`RANDOM}};
  lineBuffer_4329 = _RAND_4336[7:0];
  _RAND_4337 = {1{`RANDOM}};
  lineBuffer_4330 = _RAND_4337[7:0];
  _RAND_4338 = {1{`RANDOM}};
  lineBuffer_4331 = _RAND_4338[7:0];
  _RAND_4339 = {1{`RANDOM}};
  lineBuffer_4332 = _RAND_4339[7:0];
  _RAND_4340 = {1{`RANDOM}};
  lineBuffer_4333 = _RAND_4340[7:0];
  _RAND_4341 = {1{`RANDOM}};
  lineBuffer_4334 = _RAND_4341[7:0];
  _RAND_4342 = {1{`RANDOM}};
  lineBuffer_4335 = _RAND_4342[7:0];
  _RAND_4343 = {1{`RANDOM}};
  lineBuffer_4336 = _RAND_4343[7:0];
  _RAND_4344 = {1{`RANDOM}};
  lineBuffer_4337 = _RAND_4344[7:0];
  _RAND_4345 = {1{`RANDOM}};
  lineBuffer_4338 = _RAND_4345[7:0];
  _RAND_4346 = {1{`RANDOM}};
  lineBuffer_4339 = _RAND_4346[7:0];
  _RAND_4347 = {1{`RANDOM}};
  lineBuffer_4340 = _RAND_4347[7:0];
  _RAND_4348 = {1{`RANDOM}};
  lineBuffer_4341 = _RAND_4348[7:0];
  _RAND_4349 = {1{`RANDOM}};
  lineBuffer_4342 = _RAND_4349[7:0];
  _RAND_4350 = {1{`RANDOM}};
  lineBuffer_4343 = _RAND_4350[7:0];
  _RAND_4351 = {1{`RANDOM}};
  lineBuffer_4344 = _RAND_4351[7:0];
  _RAND_4352 = {1{`RANDOM}};
  lineBuffer_4345 = _RAND_4352[7:0];
  _RAND_4353 = {1{`RANDOM}};
  lineBuffer_4346 = _RAND_4353[7:0];
  _RAND_4354 = {1{`RANDOM}};
  lineBuffer_4347 = _RAND_4354[7:0];
  _RAND_4355 = {1{`RANDOM}};
  lineBuffer_4348 = _RAND_4355[7:0];
  _RAND_4356 = {1{`RANDOM}};
  lineBuffer_4349 = _RAND_4356[7:0];
  _RAND_4357 = {1{`RANDOM}};
  lineBuffer_4350 = _RAND_4357[7:0];
  _RAND_4358 = {1{`RANDOM}};
  lineBuffer_4351 = _RAND_4358[7:0];
  _RAND_4359 = {1{`RANDOM}};
  lineBuffer_4352 = _RAND_4359[7:0];
  _RAND_4360 = {1{`RANDOM}};
  lineBuffer_4353 = _RAND_4360[7:0];
  _RAND_4361 = {1{`RANDOM}};
  lineBuffer_4354 = _RAND_4361[7:0];
  _RAND_4362 = {1{`RANDOM}};
  lineBuffer_4355 = _RAND_4362[7:0];
  _RAND_4363 = {1{`RANDOM}};
  lineBuffer_4356 = _RAND_4363[7:0];
  _RAND_4364 = {1{`RANDOM}};
  lineBuffer_4357 = _RAND_4364[7:0];
  _RAND_4365 = {1{`RANDOM}};
  lineBuffer_4358 = _RAND_4365[7:0];
  _RAND_4366 = {1{`RANDOM}};
  lineBuffer_4359 = _RAND_4366[7:0];
  _RAND_4367 = {1{`RANDOM}};
  lineBuffer_4360 = _RAND_4367[7:0];
  _RAND_4368 = {1{`RANDOM}};
  lineBuffer_4361 = _RAND_4368[7:0];
  _RAND_4369 = {1{`RANDOM}};
  lineBuffer_4362 = _RAND_4369[7:0];
  _RAND_4370 = {1{`RANDOM}};
  lineBuffer_4363 = _RAND_4370[7:0];
  _RAND_4371 = {1{`RANDOM}};
  lineBuffer_4364 = _RAND_4371[7:0];
  _RAND_4372 = {1{`RANDOM}};
  lineBuffer_4365 = _RAND_4372[7:0];
  _RAND_4373 = {1{`RANDOM}};
  lineBuffer_4366 = _RAND_4373[7:0];
  _RAND_4374 = {1{`RANDOM}};
  lineBuffer_4367 = _RAND_4374[7:0];
  _RAND_4375 = {1{`RANDOM}};
  lineBuffer_4368 = _RAND_4375[7:0];
  _RAND_4376 = {1{`RANDOM}};
  lineBuffer_4369 = _RAND_4376[7:0];
  _RAND_4377 = {1{`RANDOM}};
  lineBuffer_4370 = _RAND_4377[7:0];
  _RAND_4378 = {1{`RANDOM}};
  lineBuffer_4371 = _RAND_4378[7:0];
  _RAND_4379 = {1{`RANDOM}};
  lineBuffer_4372 = _RAND_4379[7:0];
  _RAND_4380 = {1{`RANDOM}};
  lineBuffer_4373 = _RAND_4380[7:0];
  _RAND_4381 = {1{`RANDOM}};
  lineBuffer_4374 = _RAND_4381[7:0];
  _RAND_4382 = {1{`RANDOM}};
  lineBuffer_4375 = _RAND_4382[7:0];
  _RAND_4383 = {1{`RANDOM}};
  lineBuffer_4376 = _RAND_4383[7:0];
  _RAND_4384 = {1{`RANDOM}};
  lineBuffer_4377 = _RAND_4384[7:0];
  _RAND_4385 = {1{`RANDOM}};
  lineBuffer_4378 = _RAND_4385[7:0];
  _RAND_4386 = {1{`RANDOM}};
  lineBuffer_4379 = _RAND_4386[7:0];
  _RAND_4387 = {1{`RANDOM}};
  lineBuffer_4380 = _RAND_4387[7:0];
  _RAND_4388 = {1{`RANDOM}};
  lineBuffer_4381 = _RAND_4388[7:0];
  _RAND_4389 = {1{`RANDOM}};
  lineBuffer_4382 = _RAND_4389[7:0];
  _RAND_4390 = {1{`RANDOM}};
  lineBuffer_4383 = _RAND_4390[7:0];
  _RAND_4391 = {1{`RANDOM}};
  lineBuffer_4384 = _RAND_4391[7:0];
  _RAND_4392 = {1{`RANDOM}};
  lineBuffer_4385 = _RAND_4392[7:0];
  _RAND_4393 = {1{`RANDOM}};
  lineBuffer_4386 = _RAND_4393[7:0];
  _RAND_4394 = {1{`RANDOM}};
  lineBuffer_4387 = _RAND_4394[7:0];
  _RAND_4395 = {1{`RANDOM}};
  lineBuffer_4388 = _RAND_4395[7:0];
  _RAND_4396 = {1{`RANDOM}};
  lineBuffer_4389 = _RAND_4396[7:0];
  _RAND_4397 = {1{`RANDOM}};
  lineBuffer_4390 = _RAND_4397[7:0];
  _RAND_4398 = {1{`RANDOM}};
  lineBuffer_4391 = _RAND_4398[7:0];
  _RAND_4399 = {1{`RANDOM}};
  lineBuffer_4392 = _RAND_4399[7:0];
  _RAND_4400 = {1{`RANDOM}};
  lineBuffer_4393 = _RAND_4400[7:0];
  _RAND_4401 = {1{`RANDOM}};
  lineBuffer_4394 = _RAND_4401[7:0];
  _RAND_4402 = {1{`RANDOM}};
  lineBuffer_4395 = _RAND_4402[7:0];
  _RAND_4403 = {1{`RANDOM}};
  lineBuffer_4396 = _RAND_4403[7:0];
  _RAND_4404 = {1{`RANDOM}};
  lineBuffer_4397 = _RAND_4404[7:0];
  _RAND_4405 = {1{`RANDOM}};
  lineBuffer_4398 = _RAND_4405[7:0];
  _RAND_4406 = {1{`RANDOM}};
  lineBuffer_4399 = _RAND_4406[7:0];
  _RAND_4407 = {1{`RANDOM}};
  lineBuffer_4400 = _RAND_4407[7:0];
  _RAND_4408 = {1{`RANDOM}};
  lineBuffer_4401 = _RAND_4408[7:0];
  _RAND_4409 = {1{`RANDOM}};
  lineBuffer_4402 = _RAND_4409[7:0];
  _RAND_4410 = {1{`RANDOM}};
  lineBuffer_4403 = _RAND_4410[7:0];
  _RAND_4411 = {1{`RANDOM}};
  lineBuffer_4404 = _RAND_4411[7:0];
  _RAND_4412 = {1{`RANDOM}};
  lineBuffer_4405 = _RAND_4412[7:0];
  _RAND_4413 = {1{`RANDOM}};
  lineBuffer_4406 = _RAND_4413[7:0];
  _RAND_4414 = {1{`RANDOM}};
  lineBuffer_4407 = _RAND_4414[7:0];
  _RAND_4415 = {1{`RANDOM}};
  lineBuffer_4408 = _RAND_4415[7:0];
  _RAND_4416 = {1{`RANDOM}};
  lineBuffer_4409 = _RAND_4416[7:0];
  _RAND_4417 = {1{`RANDOM}};
  lineBuffer_4410 = _RAND_4417[7:0];
  _RAND_4418 = {1{`RANDOM}};
  lineBuffer_4411 = _RAND_4418[7:0];
  _RAND_4419 = {1{`RANDOM}};
  lineBuffer_4412 = _RAND_4419[7:0];
  _RAND_4420 = {1{`RANDOM}};
  lineBuffer_4413 = _RAND_4420[7:0];
  _RAND_4421 = {1{`RANDOM}};
  lineBuffer_4414 = _RAND_4421[7:0];
  _RAND_4422 = {1{`RANDOM}};
  lineBuffer_4415 = _RAND_4422[7:0];
  _RAND_4423 = {1{`RANDOM}};
  lineBuffer_4416 = _RAND_4423[7:0];
  _RAND_4424 = {1{`RANDOM}};
  lineBuffer_4417 = _RAND_4424[7:0];
  _RAND_4425 = {1{`RANDOM}};
  lineBuffer_4418 = _RAND_4425[7:0];
  _RAND_4426 = {1{`RANDOM}};
  lineBuffer_4419 = _RAND_4426[7:0];
  _RAND_4427 = {1{`RANDOM}};
  lineBuffer_4420 = _RAND_4427[7:0];
  _RAND_4428 = {1{`RANDOM}};
  lineBuffer_4421 = _RAND_4428[7:0];
  _RAND_4429 = {1{`RANDOM}};
  lineBuffer_4422 = _RAND_4429[7:0];
  _RAND_4430 = {1{`RANDOM}};
  lineBuffer_4423 = _RAND_4430[7:0];
  _RAND_4431 = {1{`RANDOM}};
  lineBuffer_4424 = _RAND_4431[7:0];
  _RAND_4432 = {1{`RANDOM}};
  lineBuffer_4425 = _RAND_4432[7:0];
  _RAND_4433 = {1{`RANDOM}};
  lineBuffer_4426 = _RAND_4433[7:0];
  _RAND_4434 = {1{`RANDOM}};
  lineBuffer_4427 = _RAND_4434[7:0];
  _RAND_4435 = {1{`RANDOM}};
  lineBuffer_4428 = _RAND_4435[7:0];
  _RAND_4436 = {1{`RANDOM}};
  lineBuffer_4429 = _RAND_4436[7:0];
  _RAND_4437 = {1{`RANDOM}};
  lineBuffer_4430 = _RAND_4437[7:0];
  _RAND_4438 = {1{`RANDOM}};
  lineBuffer_4431 = _RAND_4438[7:0];
  _RAND_4439 = {1{`RANDOM}};
  lineBuffer_4432 = _RAND_4439[7:0];
  _RAND_4440 = {1{`RANDOM}};
  lineBuffer_4433 = _RAND_4440[7:0];
  _RAND_4441 = {1{`RANDOM}};
  lineBuffer_4434 = _RAND_4441[7:0];
  _RAND_4442 = {1{`RANDOM}};
  lineBuffer_4435 = _RAND_4442[7:0];
  _RAND_4443 = {1{`RANDOM}};
  lineBuffer_4436 = _RAND_4443[7:0];
  _RAND_4444 = {1{`RANDOM}};
  lineBuffer_4437 = _RAND_4444[7:0];
  _RAND_4445 = {1{`RANDOM}};
  lineBuffer_4438 = _RAND_4445[7:0];
  _RAND_4446 = {1{`RANDOM}};
  lineBuffer_4439 = _RAND_4446[7:0];
  _RAND_4447 = {1{`RANDOM}};
  lineBuffer_4440 = _RAND_4447[7:0];
  _RAND_4448 = {1{`RANDOM}};
  lineBuffer_4441 = _RAND_4448[7:0];
  _RAND_4449 = {1{`RANDOM}};
  lineBuffer_4442 = _RAND_4449[7:0];
  _RAND_4450 = {1{`RANDOM}};
  lineBuffer_4443 = _RAND_4450[7:0];
  _RAND_4451 = {1{`RANDOM}};
  lineBuffer_4444 = _RAND_4451[7:0];
  _RAND_4452 = {1{`RANDOM}};
  lineBuffer_4445 = _RAND_4452[7:0];
  _RAND_4453 = {1{`RANDOM}};
  lineBuffer_4446 = _RAND_4453[7:0];
  _RAND_4454 = {1{`RANDOM}};
  lineBuffer_4447 = _RAND_4454[7:0];
  _RAND_4455 = {1{`RANDOM}};
  lineBuffer_4448 = _RAND_4455[7:0];
  _RAND_4456 = {1{`RANDOM}};
  lineBuffer_4449 = _RAND_4456[7:0];
  _RAND_4457 = {1{`RANDOM}};
  lineBuffer_4450 = _RAND_4457[7:0];
  _RAND_4458 = {1{`RANDOM}};
  lineBuffer_4451 = _RAND_4458[7:0];
  _RAND_4459 = {1{`RANDOM}};
  lineBuffer_4452 = _RAND_4459[7:0];
  _RAND_4460 = {1{`RANDOM}};
  lineBuffer_4453 = _RAND_4460[7:0];
  _RAND_4461 = {1{`RANDOM}};
  lineBuffer_4454 = _RAND_4461[7:0];
  _RAND_4462 = {1{`RANDOM}};
  lineBuffer_4455 = _RAND_4462[7:0];
  _RAND_4463 = {1{`RANDOM}};
  lineBuffer_4456 = _RAND_4463[7:0];
  _RAND_4464 = {1{`RANDOM}};
  lineBuffer_4457 = _RAND_4464[7:0];
  _RAND_4465 = {1{`RANDOM}};
  lineBuffer_4458 = _RAND_4465[7:0];
  _RAND_4466 = {1{`RANDOM}};
  lineBuffer_4459 = _RAND_4466[7:0];
  _RAND_4467 = {1{`RANDOM}};
  lineBuffer_4460 = _RAND_4467[7:0];
  _RAND_4468 = {1{`RANDOM}};
  lineBuffer_4461 = _RAND_4468[7:0];
  _RAND_4469 = {1{`RANDOM}};
  lineBuffer_4462 = _RAND_4469[7:0];
  _RAND_4470 = {1{`RANDOM}};
  lineBuffer_4463 = _RAND_4470[7:0];
  _RAND_4471 = {1{`RANDOM}};
  lineBuffer_4464 = _RAND_4471[7:0];
  _RAND_4472 = {1{`RANDOM}};
  lineBuffer_4465 = _RAND_4472[7:0];
  _RAND_4473 = {1{`RANDOM}};
  lineBuffer_4466 = _RAND_4473[7:0];
  _RAND_4474 = {1{`RANDOM}};
  lineBuffer_4467 = _RAND_4474[7:0];
  _RAND_4475 = {1{`RANDOM}};
  lineBuffer_4468 = _RAND_4475[7:0];
  _RAND_4476 = {1{`RANDOM}};
  lineBuffer_4469 = _RAND_4476[7:0];
  _RAND_4477 = {1{`RANDOM}};
  lineBuffer_4470 = _RAND_4477[7:0];
  _RAND_4478 = {1{`RANDOM}};
  lineBuffer_4471 = _RAND_4478[7:0];
  _RAND_4479 = {1{`RANDOM}};
  lineBuffer_4472 = _RAND_4479[7:0];
  _RAND_4480 = {1{`RANDOM}};
  lineBuffer_4473 = _RAND_4480[7:0];
  _RAND_4481 = {1{`RANDOM}};
  lineBuffer_4474 = _RAND_4481[7:0];
  _RAND_4482 = {1{`RANDOM}};
  lineBuffer_4475 = _RAND_4482[7:0];
  _RAND_4483 = {1{`RANDOM}};
  lineBuffer_4476 = _RAND_4483[7:0];
  _RAND_4484 = {1{`RANDOM}};
  lineBuffer_4477 = _RAND_4484[7:0];
  _RAND_4485 = {1{`RANDOM}};
  lineBuffer_4478 = _RAND_4485[7:0];
  _RAND_4486 = {1{`RANDOM}};
  lineBuffer_4479 = _RAND_4486[7:0];
  _RAND_4487 = {1{`RANDOM}};
  lineBuffer_4480 = _RAND_4487[7:0];
  _RAND_4488 = {1{`RANDOM}};
  lineBuffer_4481 = _RAND_4488[7:0];
  _RAND_4489 = {1{`RANDOM}};
  lineBuffer_4482 = _RAND_4489[7:0];
  _RAND_4490 = {1{`RANDOM}};
  lineBuffer_4483 = _RAND_4490[7:0];
  _RAND_4491 = {1{`RANDOM}};
  lineBuffer_4484 = _RAND_4491[7:0];
  _RAND_4492 = {1{`RANDOM}};
  lineBuffer_4485 = _RAND_4492[7:0];
  _RAND_4493 = {1{`RANDOM}};
  lineBuffer_4486 = _RAND_4493[7:0];
  _RAND_4494 = {1{`RANDOM}};
  lineBuffer_4487 = _RAND_4494[7:0];
  _RAND_4495 = {1{`RANDOM}};
  lineBuffer_4488 = _RAND_4495[7:0];
  _RAND_4496 = {1{`RANDOM}};
  lineBuffer_4489 = _RAND_4496[7:0];
  _RAND_4497 = {1{`RANDOM}};
  lineBuffer_4490 = _RAND_4497[7:0];
  _RAND_4498 = {1{`RANDOM}};
  lineBuffer_4491 = _RAND_4498[7:0];
  _RAND_4499 = {1{`RANDOM}};
  lineBuffer_4492 = _RAND_4499[7:0];
  _RAND_4500 = {1{`RANDOM}};
  lineBuffer_4493 = _RAND_4500[7:0];
  _RAND_4501 = {1{`RANDOM}};
  lineBuffer_4494 = _RAND_4501[7:0];
  _RAND_4502 = {1{`RANDOM}};
  lineBuffer_4495 = _RAND_4502[7:0];
  _RAND_4503 = {1{`RANDOM}};
  lineBuffer_4496 = _RAND_4503[7:0];
  _RAND_4504 = {1{`RANDOM}};
  lineBuffer_4497 = _RAND_4504[7:0];
  _RAND_4505 = {1{`RANDOM}};
  lineBuffer_4498 = _RAND_4505[7:0];
  _RAND_4506 = {1{`RANDOM}};
  lineBuffer_4499 = _RAND_4506[7:0];
  _RAND_4507 = {1{`RANDOM}};
  lineBuffer_4500 = _RAND_4507[7:0];
  _RAND_4508 = {1{`RANDOM}};
  lineBuffer_4501 = _RAND_4508[7:0];
  _RAND_4509 = {1{`RANDOM}};
  lineBuffer_4502 = _RAND_4509[7:0];
  _RAND_4510 = {1{`RANDOM}};
  lineBuffer_4503 = _RAND_4510[7:0];
  _RAND_4511 = {1{`RANDOM}};
  lineBuffer_4504 = _RAND_4511[7:0];
  _RAND_4512 = {1{`RANDOM}};
  lineBuffer_4505 = _RAND_4512[7:0];
  _RAND_4513 = {1{`RANDOM}};
  lineBuffer_4506 = _RAND_4513[7:0];
  _RAND_4514 = {1{`RANDOM}};
  lineBuffer_4507 = _RAND_4514[7:0];
  _RAND_4515 = {1{`RANDOM}};
  lineBuffer_4508 = _RAND_4515[7:0];
  _RAND_4516 = {1{`RANDOM}};
  lineBuffer_4509 = _RAND_4516[7:0];
  _RAND_4517 = {1{`RANDOM}};
  lineBuffer_4510 = _RAND_4517[7:0];
  _RAND_4518 = {1{`RANDOM}};
  lineBuffer_4511 = _RAND_4518[7:0];
  _RAND_4519 = {1{`RANDOM}};
  lineBuffer_4512 = _RAND_4519[7:0];
  _RAND_4520 = {1{`RANDOM}};
  lineBuffer_4513 = _RAND_4520[7:0];
  _RAND_4521 = {1{`RANDOM}};
  lineBuffer_4514 = _RAND_4521[7:0];
  _RAND_4522 = {1{`RANDOM}};
  lineBuffer_4515 = _RAND_4522[7:0];
  _RAND_4523 = {1{`RANDOM}};
  lineBuffer_4516 = _RAND_4523[7:0];
  _RAND_4524 = {1{`RANDOM}};
  lineBuffer_4517 = _RAND_4524[7:0];
  _RAND_4525 = {1{`RANDOM}};
  lineBuffer_4518 = _RAND_4525[7:0];
  _RAND_4526 = {1{`RANDOM}};
  lineBuffer_4519 = _RAND_4526[7:0];
  _RAND_4527 = {1{`RANDOM}};
  lineBuffer_4520 = _RAND_4527[7:0];
  _RAND_4528 = {1{`RANDOM}};
  lineBuffer_4521 = _RAND_4528[7:0];
  _RAND_4529 = {1{`RANDOM}};
  lineBuffer_4522 = _RAND_4529[7:0];
  _RAND_4530 = {1{`RANDOM}};
  lineBuffer_4523 = _RAND_4530[7:0];
  _RAND_4531 = {1{`RANDOM}};
  lineBuffer_4524 = _RAND_4531[7:0];
  _RAND_4532 = {1{`RANDOM}};
  lineBuffer_4525 = _RAND_4532[7:0];
  _RAND_4533 = {1{`RANDOM}};
  lineBuffer_4526 = _RAND_4533[7:0];
  _RAND_4534 = {1{`RANDOM}};
  lineBuffer_4527 = _RAND_4534[7:0];
  _RAND_4535 = {1{`RANDOM}};
  lineBuffer_4528 = _RAND_4535[7:0];
  _RAND_4536 = {1{`RANDOM}};
  lineBuffer_4529 = _RAND_4536[7:0];
  _RAND_4537 = {1{`RANDOM}};
  lineBuffer_4530 = _RAND_4537[7:0];
  _RAND_4538 = {1{`RANDOM}};
  lineBuffer_4531 = _RAND_4538[7:0];
  _RAND_4539 = {1{`RANDOM}};
  lineBuffer_4532 = _RAND_4539[7:0];
  _RAND_4540 = {1{`RANDOM}};
  lineBuffer_4533 = _RAND_4540[7:0];
  _RAND_4541 = {1{`RANDOM}};
  lineBuffer_4534 = _RAND_4541[7:0];
  _RAND_4542 = {1{`RANDOM}};
  lineBuffer_4535 = _RAND_4542[7:0];
  _RAND_4543 = {1{`RANDOM}};
  lineBuffer_4536 = _RAND_4543[7:0];
  _RAND_4544 = {1{`RANDOM}};
  lineBuffer_4537 = _RAND_4544[7:0];
  _RAND_4545 = {1{`RANDOM}};
  lineBuffer_4538 = _RAND_4545[7:0];
  _RAND_4546 = {1{`RANDOM}};
  lineBuffer_4539 = _RAND_4546[7:0];
  _RAND_4547 = {1{`RANDOM}};
  lineBuffer_4540 = _RAND_4547[7:0];
  _RAND_4548 = {1{`RANDOM}};
  lineBuffer_4541 = _RAND_4548[7:0];
  _RAND_4549 = {1{`RANDOM}};
  lineBuffer_4542 = _RAND_4549[7:0];
  _RAND_4550 = {1{`RANDOM}};
  lineBuffer_4543 = _RAND_4550[7:0];
  _RAND_4551 = {1{`RANDOM}};
  lineBuffer_4544 = _RAND_4551[7:0];
  _RAND_4552 = {1{`RANDOM}};
  lineBuffer_4545 = _RAND_4552[7:0];
  _RAND_4553 = {1{`RANDOM}};
  lineBuffer_4546 = _RAND_4553[7:0];
  _RAND_4554 = {1{`RANDOM}};
  lineBuffer_4547 = _RAND_4554[7:0];
  _RAND_4555 = {1{`RANDOM}};
  lineBuffer_4548 = _RAND_4555[7:0];
  _RAND_4556 = {1{`RANDOM}};
  lineBuffer_4549 = _RAND_4556[7:0];
  _RAND_4557 = {1{`RANDOM}};
  lineBuffer_4550 = _RAND_4557[7:0];
  _RAND_4558 = {1{`RANDOM}};
  lineBuffer_4551 = _RAND_4558[7:0];
  _RAND_4559 = {1{`RANDOM}};
  lineBuffer_4552 = _RAND_4559[7:0];
  _RAND_4560 = {1{`RANDOM}};
  lineBuffer_4553 = _RAND_4560[7:0];
  _RAND_4561 = {1{`RANDOM}};
  lineBuffer_4554 = _RAND_4561[7:0];
  _RAND_4562 = {1{`RANDOM}};
  lineBuffer_4555 = _RAND_4562[7:0];
  _RAND_4563 = {1{`RANDOM}};
  lineBuffer_4556 = _RAND_4563[7:0];
  _RAND_4564 = {1{`RANDOM}};
  lineBuffer_4557 = _RAND_4564[7:0];
  _RAND_4565 = {1{`RANDOM}};
  lineBuffer_4558 = _RAND_4565[7:0];
  _RAND_4566 = {1{`RANDOM}};
  lineBuffer_4559 = _RAND_4566[7:0];
  _RAND_4567 = {1{`RANDOM}};
  lineBuffer_4560 = _RAND_4567[7:0];
  _RAND_4568 = {1{`RANDOM}};
  lineBuffer_4561 = _RAND_4568[7:0];
  _RAND_4569 = {1{`RANDOM}};
  lineBuffer_4562 = _RAND_4569[7:0];
  _RAND_4570 = {1{`RANDOM}};
  lineBuffer_4563 = _RAND_4570[7:0];
  _RAND_4571 = {1{`RANDOM}};
  lineBuffer_4564 = _RAND_4571[7:0];
  _RAND_4572 = {1{`RANDOM}};
  lineBuffer_4565 = _RAND_4572[7:0];
  _RAND_4573 = {1{`RANDOM}};
  lineBuffer_4566 = _RAND_4573[7:0];
  _RAND_4574 = {1{`RANDOM}};
  lineBuffer_4567 = _RAND_4574[7:0];
  _RAND_4575 = {1{`RANDOM}};
  lineBuffer_4568 = _RAND_4575[7:0];
  _RAND_4576 = {1{`RANDOM}};
  lineBuffer_4569 = _RAND_4576[7:0];
  _RAND_4577 = {1{`RANDOM}};
  lineBuffer_4570 = _RAND_4577[7:0];
  _RAND_4578 = {1{`RANDOM}};
  lineBuffer_4571 = _RAND_4578[7:0];
  _RAND_4579 = {1{`RANDOM}};
  lineBuffer_4572 = _RAND_4579[7:0];
  _RAND_4580 = {1{`RANDOM}};
  lineBuffer_4573 = _RAND_4580[7:0];
  _RAND_4581 = {1{`RANDOM}};
  lineBuffer_4574 = _RAND_4581[7:0];
  _RAND_4582 = {1{`RANDOM}};
  lineBuffer_4575 = _RAND_4582[7:0];
  _RAND_4583 = {1{`RANDOM}};
  lineBuffer_4576 = _RAND_4583[7:0];
  _RAND_4584 = {1{`RANDOM}};
  lineBuffer_4577 = _RAND_4584[7:0];
  _RAND_4585 = {1{`RANDOM}};
  lineBuffer_4578 = _RAND_4585[7:0];
  _RAND_4586 = {1{`RANDOM}};
  lineBuffer_4579 = _RAND_4586[7:0];
  _RAND_4587 = {1{`RANDOM}};
  lineBuffer_4580 = _RAND_4587[7:0];
  _RAND_4588 = {1{`RANDOM}};
  lineBuffer_4581 = _RAND_4588[7:0];
  _RAND_4589 = {1{`RANDOM}};
  lineBuffer_4582 = _RAND_4589[7:0];
  _RAND_4590 = {1{`RANDOM}};
  lineBuffer_4583 = _RAND_4590[7:0];
  _RAND_4591 = {1{`RANDOM}};
  lineBuffer_4584 = _RAND_4591[7:0];
  _RAND_4592 = {1{`RANDOM}};
  lineBuffer_4585 = _RAND_4592[7:0];
  _RAND_4593 = {1{`RANDOM}};
  lineBuffer_4586 = _RAND_4593[7:0];
  _RAND_4594 = {1{`RANDOM}};
  lineBuffer_4587 = _RAND_4594[7:0];
  _RAND_4595 = {1{`RANDOM}};
  lineBuffer_4588 = _RAND_4595[7:0];
  _RAND_4596 = {1{`RANDOM}};
  lineBuffer_4589 = _RAND_4596[7:0];
  _RAND_4597 = {1{`RANDOM}};
  lineBuffer_4590 = _RAND_4597[7:0];
  _RAND_4598 = {1{`RANDOM}};
  lineBuffer_4591 = _RAND_4598[7:0];
  _RAND_4599 = {1{`RANDOM}};
  lineBuffer_4592 = _RAND_4599[7:0];
  _RAND_4600 = {1{`RANDOM}};
  lineBuffer_4593 = _RAND_4600[7:0];
  _RAND_4601 = {1{`RANDOM}};
  lineBuffer_4594 = _RAND_4601[7:0];
  _RAND_4602 = {1{`RANDOM}};
  lineBuffer_4595 = _RAND_4602[7:0];
  _RAND_4603 = {1{`RANDOM}};
  lineBuffer_4596 = _RAND_4603[7:0];
  _RAND_4604 = {1{`RANDOM}};
  lineBuffer_4597 = _RAND_4604[7:0];
  _RAND_4605 = {1{`RANDOM}};
  lineBuffer_4598 = _RAND_4605[7:0];
  _RAND_4606 = {1{`RANDOM}};
  lineBuffer_4599 = _RAND_4606[7:0];
  _RAND_4607 = {1{`RANDOM}};
  lineBuffer_4600 = _RAND_4607[7:0];
  _RAND_4608 = {1{`RANDOM}};
  lineBuffer_4601 = _RAND_4608[7:0];
  _RAND_4609 = {1{`RANDOM}};
  lineBuffer_4602 = _RAND_4609[7:0];
  _RAND_4610 = {1{`RANDOM}};
  lineBuffer_4603 = _RAND_4610[7:0];
  _RAND_4611 = {1{`RANDOM}};
  lineBuffer_4604 = _RAND_4611[7:0];
  _RAND_4612 = {1{`RANDOM}};
  lineBuffer_4605 = _RAND_4612[7:0];
  _RAND_4613 = {1{`RANDOM}};
  lineBuffer_4606 = _RAND_4613[7:0];
  _RAND_4614 = {1{`RANDOM}};
  lineBuffer_4607 = _RAND_4614[7:0];
  _RAND_4615 = {1{`RANDOM}};
  lineBuffer_4608 = _RAND_4615[7:0];
  _RAND_4616 = {1{`RANDOM}};
  lineBuffer_4609 = _RAND_4616[7:0];
  _RAND_4617 = {1{`RANDOM}};
  lineBuffer_4610 = _RAND_4617[7:0];
  _RAND_4618 = {1{`RANDOM}};
  lineBuffer_4611 = _RAND_4618[7:0];
  _RAND_4619 = {1{`RANDOM}};
  lineBuffer_4612 = _RAND_4619[7:0];
  _RAND_4620 = {1{`RANDOM}};
  lineBuffer_4613 = _RAND_4620[7:0];
  _RAND_4621 = {1{`RANDOM}};
  lineBuffer_4614 = _RAND_4621[7:0];
  _RAND_4622 = {1{`RANDOM}};
  lineBuffer_4615 = _RAND_4622[7:0];
  _RAND_4623 = {1{`RANDOM}};
  lineBuffer_4616 = _RAND_4623[7:0];
  _RAND_4624 = {1{`RANDOM}};
  lineBuffer_4617 = _RAND_4624[7:0];
  _RAND_4625 = {1{`RANDOM}};
  lineBuffer_4618 = _RAND_4625[7:0];
  _RAND_4626 = {1{`RANDOM}};
  lineBuffer_4619 = _RAND_4626[7:0];
  _RAND_4627 = {1{`RANDOM}};
  lineBuffer_4620 = _RAND_4627[7:0];
  _RAND_4628 = {1{`RANDOM}};
  lineBuffer_4621 = _RAND_4628[7:0];
  _RAND_4629 = {1{`RANDOM}};
  lineBuffer_4622 = _RAND_4629[7:0];
  _RAND_4630 = {1{`RANDOM}};
  lineBuffer_4623 = _RAND_4630[7:0];
  _RAND_4631 = {1{`RANDOM}};
  lineBuffer_4624 = _RAND_4631[7:0];
  _RAND_4632 = {1{`RANDOM}};
  lineBuffer_4625 = _RAND_4632[7:0];
  _RAND_4633 = {1{`RANDOM}};
  lineBuffer_4626 = _RAND_4633[7:0];
  _RAND_4634 = {1{`RANDOM}};
  lineBuffer_4627 = _RAND_4634[7:0];
  _RAND_4635 = {1{`RANDOM}};
  lineBuffer_4628 = _RAND_4635[7:0];
  _RAND_4636 = {1{`RANDOM}};
  lineBuffer_4629 = _RAND_4636[7:0];
  _RAND_4637 = {1{`RANDOM}};
  lineBuffer_4630 = _RAND_4637[7:0];
  _RAND_4638 = {1{`RANDOM}};
  lineBuffer_4631 = _RAND_4638[7:0];
  _RAND_4639 = {1{`RANDOM}};
  lineBuffer_4632 = _RAND_4639[7:0];
  _RAND_4640 = {1{`RANDOM}};
  lineBuffer_4633 = _RAND_4640[7:0];
  _RAND_4641 = {1{`RANDOM}};
  lineBuffer_4634 = _RAND_4641[7:0];
  _RAND_4642 = {1{`RANDOM}};
  lineBuffer_4635 = _RAND_4642[7:0];
  _RAND_4643 = {1{`RANDOM}};
  lineBuffer_4636 = _RAND_4643[7:0];
  _RAND_4644 = {1{`RANDOM}};
  lineBuffer_4637 = _RAND_4644[7:0];
  _RAND_4645 = {1{`RANDOM}};
  lineBuffer_4638 = _RAND_4645[7:0];
  _RAND_4646 = {1{`RANDOM}};
  lineBuffer_4639 = _RAND_4646[7:0];
  _RAND_4647 = {1{`RANDOM}};
  lineBuffer_4640 = _RAND_4647[7:0];
  _RAND_4648 = {1{`RANDOM}};
  lineBuffer_4641 = _RAND_4648[7:0];
  _RAND_4649 = {1{`RANDOM}};
  lineBuffer_4642 = _RAND_4649[7:0];
  _RAND_4650 = {1{`RANDOM}};
  lineBuffer_4643 = _RAND_4650[7:0];
  _RAND_4651 = {1{`RANDOM}};
  lineBuffer_4644 = _RAND_4651[7:0];
  _RAND_4652 = {1{`RANDOM}};
  lineBuffer_4645 = _RAND_4652[7:0];
  _RAND_4653 = {1{`RANDOM}};
  lineBuffer_4646 = _RAND_4653[7:0];
  _RAND_4654 = {1{`RANDOM}};
  lineBuffer_4647 = _RAND_4654[7:0];
  _RAND_4655 = {1{`RANDOM}};
  lineBuffer_4648 = _RAND_4655[7:0];
  _RAND_4656 = {1{`RANDOM}};
  lineBuffer_4649 = _RAND_4656[7:0];
  _RAND_4657 = {1{`RANDOM}};
  lineBuffer_4650 = _RAND_4657[7:0];
  _RAND_4658 = {1{`RANDOM}};
  lineBuffer_4651 = _RAND_4658[7:0];
  _RAND_4659 = {1{`RANDOM}};
  lineBuffer_4652 = _RAND_4659[7:0];
  _RAND_4660 = {1{`RANDOM}};
  lineBuffer_4653 = _RAND_4660[7:0];
  _RAND_4661 = {1{`RANDOM}};
  lineBuffer_4654 = _RAND_4661[7:0];
  _RAND_4662 = {1{`RANDOM}};
  lineBuffer_4655 = _RAND_4662[7:0];
  _RAND_4663 = {1{`RANDOM}};
  lineBuffer_4656 = _RAND_4663[7:0];
  _RAND_4664 = {1{`RANDOM}};
  lineBuffer_4657 = _RAND_4664[7:0];
  _RAND_4665 = {1{`RANDOM}};
  lineBuffer_4658 = _RAND_4665[7:0];
  _RAND_4666 = {1{`RANDOM}};
  lineBuffer_4659 = _RAND_4666[7:0];
  _RAND_4667 = {1{`RANDOM}};
  lineBuffer_4660 = _RAND_4667[7:0];
  _RAND_4668 = {1{`RANDOM}};
  lineBuffer_4661 = _RAND_4668[7:0];
  _RAND_4669 = {1{`RANDOM}};
  lineBuffer_4662 = _RAND_4669[7:0];
  _RAND_4670 = {1{`RANDOM}};
  lineBuffer_4663 = _RAND_4670[7:0];
  _RAND_4671 = {1{`RANDOM}};
  lineBuffer_4664 = _RAND_4671[7:0];
  _RAND_4672 = {1{`RANDOM}};
  lineBuffer_4665 = _RAND_4672[7:0];
  _RAND_4673 = {1{`RANDOM}};
  lineBuffer_4666 = _RAND_4673[7:0];
  _RAND_4674 = {1{`RANDOM}};
  lineBuffer_4667 = _RAND_4674[7:0];
  _RAND_4675 = {1{`RANDOM}};
  lineBuffer_4668 = _RAND_4675[7:0];
  _RAND_4676 = {1{`RANDOM}};
  lineBuffer_4669 = _RAND_4676[7:0];
  _RAND_4677 = {1{`RANDOM}};
  lineBuffer_4670 = _RAND_4677[7:0];
  _RAND_4678 = {1{`RANDOM}};
  lineBuffer_4671 = _RAND_4678[7:0];
  _RAND_4679 = {1{`RANDOM}};
  lineBuffer_4672 = _RAND_4679[7:0];
  _RAND_4680 = {1{`RANDOM}};
  lineBuffer_4673 = _RAND_4680[7:0];
  _RAND_4681 = {1{`RANDOM}};
  lineBuffer_4674 = _RAND_4681[7:0];
  _RAND_4682 = {1{`RANDOM}};
  lineBuffer_4675 = _RAND_4682[7:0];
  _RAND_4683 = {1{`RANDOM}};
  lineBuffer_4676 = _RAND_4683[7:0];
  _RAND_4684 = {1{`RANDOM}};
  lineBuffer_4677 = _RAND_4684[7:0];
  _RAND_4685 = {1{`RANDOM}};
  lineBuffer_4678 = _RAND_4685[7:0];
  _RAND_4686 = {1{`RANDOM}};
  lineBuffer_4679 = _RAND_4686[7:0];
  _RAND_4687 = {1{`RANDOM}};
  lineBuffer_4680 = _RAND_4687[7:0];
  _RAND_4688 = {1{`RANDOM}};
  lineBuffer_4681 = _RAND_4688[7:0];
  _RAND_4689 = {1{`RANDOM}};
  lineBuffer_4682 = _RAND_4689[7:0];
  _RAND_4690 = {1{`RANDOM}};
  lineBuffer_4683 = _RAND_4690[7:0];
  _RAND_4691 = {1{`RANDOM}};
  lineBuffer_4684 = _RAND_4691[7:0];
  _RAND_4692 = {1{`RANDOM}};
  lineBuffer_4685 = _RAND_4692[7:0];
  _RAND_4693 = {1{`RANDOM}};
  lineBuffer_4686 = _RAND_4693[7:0];
  _RAND_4694 = {1{`RANDOM}};
  lineBuffer_4687 = _RAND_4694[7:0];
  _RAND_4695 = {1{`RANDOM}};
  lineBuffer_4688 = _RAND_4695[7:0];
  _RAND_4696 = {1{`RANDOM}};
  lineBuffer_4689 = _RAND_4696[7:0];
  _RAND_4697 = {1{`RANDOM}};
  lineBuffer_4690 = _RAND_4697[7:0];
  _RAND_4698 = {1{`RANDOM}};
  lineBuffer_4691 = _RAND_4698[7:0];
  _RAND_4699 = {1{`RANDOM}};
  lineBuffer_4692 = _RAND_4699[7:0];
  _RAND_4700 = {1{`RANDOM}};
  lineBuffer_4693 = _RAND_4700[7:0];
  _RAND_4701 = {1{`RANDOM}};
  lineBuffer_4694 = _RAND_4701[7:0];
  _RAND_4702 = {1{`RANDOM}};
  lineBuffer_4695 = _RAND_4702[7:0];
  _RAND_4703 = {1{`RANDOM}};
  lineBuffer_4696 = _RAND_4703[7:0];
  _RAND_4704 = {1{`RANDOM}};
  lineBuffer_4697 = _RAND_4704[7:0];
  _RAND_4705 = {1{`RANDOM}};
  lineBuffer_4698 = _RAND_4705[7:0];
  _RAND_4706 = {1{`RANDOM}};
  lineBuffer_4699 = _RAND_4706[7:0];
  _RAND_4707 = {1{`RANDOM}};
  lineBuffer_4700 = _RAND_4707[7:0];
  _RAND_4708 = {1{`RANDOM}};
  lineBuffer_4701 = _RAND_4708[7:0];
  _RAND_4709 = {1{`RANDOM}};
  lineBuffer_4702 = _RAND_4709[7:0];
  _RAND_4710 = {1{`RANDOM}};
  lineBuffer_4703 = _RAND_4710[7:0];
  _RAND_4711 = {1{`RANDOM}};
  lineBuffer_4704 = _RAND_4711[7:0];
  _RAND_4712 = {1{`RANDOM}};
  lineBuffer_4705 = _RAND_4712[7:0];
  _RAND_4713 = {1{`RANDOM}};
  lineBuffer_4706 = _RAND_4713[7:0];
  _RAND_4714 = {1{`RANDOM}};
  lineBuffer_4707 = _RAND_4714[7:0];
  _RAND_4715 = {1{`RANDOM}};
  lineBuffer_4708 = _RAND_4715[7:0];
  _RAND_4716 = {1{`RANDOM}};
  lineBuffer_4709 = _RAND_4716[7:0];
  _RAND_4717 = {1{`RANDOM}};
  lineBuffer_4710 = _RAND_4717[7:0];
  _RAND_4718 = {1{`RANDOM}};
  lineBuffer_4711 = _RAND_4718[7:0];
  _RAND_4719 = {1{`RANDOM}};
  lineBuffer_4712 = _RAND_4719[7:0];
  _RAND_4720 = {1{`RANDOM}};
  lineBuffer_4713 = _RAND_4720[7:0];
  _RAND_4721 = {1{`RANDOM}};
  lineBuffer_4714 = _RAND_4721[7:0];
  _RAND_4722 = {1{`RANDOM}};
  lineBuffer_4715 = _RAND_4722[7:0];
  _RAND_4723 = {1{`RANDOM}};
  lineBuffer_4716 = _RAND_4723[7:0];
  _RAND_4724 = {1{`RANDOM}};
  lineBuffer_4717 = _RAND_4724[7:0];
  _RAND_4725 = {1{`RANDOM}};
  lineBuffer_4718 = _RAND_4725[7:0];
  _RAND_4726 = {1{`RANDOM}};
  lineBuffer_4719 = _RAND_4726[7:0];
  _RAND_4727 = {1{`RANDOM}};
  lineBuffer_4720 = _RAND_4727[7:0];
  _RAND_4728 = {1{`RANDOM}};
  lineBuffer_4721 = _RAND_4728[7:0];
  _RAND_4729 = {1{`RANDOM}};
  lineBuffer_4722 = _RAND_4729[7:0];
  _RAND_4730 = {1{`RANDOM}};
  lineBuffer_4723 = _RAND_4730[7:0];
  _RAND_4731 = {1{`RANDOM}};
  lineBuffer_4724 = _RAND_4731[7:0];
  _RAND_4732 = {1{`RANDOM}};
  lineBuffer_4725 = _RAND_4732[7:0];
  _RAND_4733 = {1{`RANDOM}};
  lineBuffer_4726 = _RAND_4733[7:0];
  _RAND_4734 = {1{`RANDOM}};
  lineBuffer_4727 = _RAND_4734[7:0];
  _RAND_4735 = {1{`RANDOM}};
  lineBuffer_4728 = _RAND_4735[7:0];
  _RAND_4736 = {1{`RANDOM}};
  lineBuffer_4729 = _RAND_4736[7:0];
  _RAND_4737 = {1{`RANDOM}};
  lineBuffer_4730 = _RAND_4737[7:0];
  _RAND_4738 = {1{`RANDOM}};
  lineBuffer_4731 = _RAND_4738[7:0];
  _RAND_4739 = {1{`RANDOM}};
  lineBuffer_4732 = _RAND_4739[7:0];
  _RAND_4740 = {1{`RANDOM}};
  lineBuffer_4733 = _RAND_4740[7:0];
  _RAND_4741 = {1{`RANDOM}};
  lineBuffer_4734 = _RAND_4741[7:0];
  _RAND_4742 = {1{`RANDOM}};
  lineBuffer_4735 = _RAND_4742[7:0];
  _RAND_4743 = {1{`RANDOM}};
  lineBuffer_4736 = _RAND_4743[7:0];
  _RAND_4744 = {1{`RANDOM}};
  lineBuffer_4737 = _RAND_4744[7:0];
  _RAND_4745 = {1{`RANDOM}};
  lineBuffer_4738 = _RAND_4745[7:0];
  _RAND_4746 = {1{`RANDOM}};
  lineBuffer_4739 = _RAND_4746[7:0];
  _RAND_4747 = {1{`RANDOM}};
  lineBuffer_4740 = _RAND_4747[7:0];
  _RAND_4748 = {1{`RANDOM}};
  lineBuffer_4741 = _RAND_4748[7:0];
  _RAND_4749 = {1{`RANDOM}};
  lineBuffer_4742 = _RAND_4749[7:0];
  _RAND_4750 = {1{`RANDOM}};
  lineBuffer_4743 = _RAND_4750[7:0];
  _RAND_4751 = {1{`RANDOM}};
  lineBuffer_4744 = _RAND_4751[7:0];
  _RAND_4752 = {1{`RANDOM}};
  lineBuffer_4745 = _RAND_4752[7:0];
  _RAND_4753 = {1{`RANDOM}};
  lineBuffer_4746 = _RAND_4753[7:0];
  _RAND_4754 = {1{`RANDOM}};
  lineBuffer_4747 = _RAND_4754[7:0];
  _RAND_4755 = {1{`RANDOM}};
  lineBuffer_4748 = _RAND_4755[7:0];
  _RAND_4756 = {1{`RANDOM}};
  lineBuffer_4749 = _RAND_4756[7:0];
  _RAND_4757 = {1{`RANDOM}};
  lineBuffer_4750 = _RAND_4757[7:0];
  _RAND_4758 = {1{`RANDOM}};
  lineBuffer_4751 = _RAND_4758[7:0];
  _RAND_4759 = {1{`RANDOM}};
  lineBuffer_4752 = _RAND_4759[7:0];
  _RAND_4760 = {1{`RANDOM}};
  lineBuffer_4753 = _RAND_4760[7:0];
  _RAND_4761 = {1{`RANDOM}};
  lineBuffer_4754 = _RAND_4761[7:0];
  _RAND_4762 = {1{`RANDOM}};
  lineBuffer_4755 = _RAND_4762[7:0];
  _RAND_4763 = {1{`RANDOM}};
  lineBuffer_4756 = _RAND_4763[7:0];
  _RAND_4764 = {1{`RANDOM}};
  lineBuffer_4757 = _RAND_4764[7:0];
  _RAND_4765 = {1{`RANDOM}};
  lineBuffer_4758 = _RAND_4765[7:0];
  _RAND_4766 = {1{`RANDOM}};
  lineBuffer_4759 = _RAND_4766[7:0];
  _RAND_4767 = {1{`RANDOM}};
  lineBuffer_4760 = _RAND_4767[7:0];
  _RAND_4768 = {1{`RANDOM}};
  lineBuffer_4761 = _RAND_4768[7:0];
  _RAND_4769 = {1{`RANDOM}};
  lineBuffer_4762 = _RAND_4769[7:0];
  _RAND_4770 = {1{`RANDOM}};
  lineBuffer_4763 = _RAND_4770[7:0];
  _RAND_4771 = {1{`RANDOM}};
  lineBuffer_4764 = _RAND_4771[7:0];
  _RAND_4772 = {1{`RANDOM}};
  lineBuffer_4765 = _RAND_4772[7:0];
  _RAND_4773 = {1{`RANDOM}};
  lineBuffer_4766 = _RAND_4773[7:0];
  _RAND_4774 = {1{`RANDOM}};
  lineBuffer_4767 = _RAND_4774[7:0];
  _RAND_4775 = {1{`RANDOM}};
  lineBuffer_4768 = _RAND_4775[7:0];
  _RAND_4776 = {1{`RANDOM}};
  lineBuffer_4769 = _RAND_4776[7:0];
  _RAND_4777 = {1{`RANDOM}};
  lineBuffer_4770 = _RAND_4777[7:0];
  _RAND_4778 = {1{`RANDOM}};
  lineBuffer_4771 = _RAND_4778[7:0];
  _RAND_4779 = {1{`RANDOM}};
  lineBuffer_4772 = _RAND_4779[7:0];
  _RAND_4780 = {1{`RANDOM}};
  lineBuffer_4773 = _RAND_4780[7:0];
  _RAND_4781 = {1{`RANDOM}};
  lineBuffer_4774 = _RAND_4781[7:0];
  _RAND_4782 = {1{`RANDOM}};
  lineBuffer_4775 = _RAND_4782[7:0];
  _RAND_4783 = {1{`RANDOM}};
  lineBuffer_4776 = _RAND_4783[7:0];
  _RAND_4784 = {1{`RANDOM}};
  lineBuffer_4777 = _RAND_4784[7:0];
  _RAND_4785 = {1{`RANDOM}};
  lineBuffer_4778 = _RAND_4785[7:0];
  _RAND_4786 = {1{`RANDOM}};
  lineBuffer_4779 = _RAND_4786[7:0];
  _RAND_4787 = {1{`RANDOM}};
  lineBuffer_4780 = _RAND_4787[7:0];
  _RAND_4788 = {1{`RANDOM}};
  lineBuffer_4781 = _RAND_4788[7:0];
  _RAND_4789 = {1{`RANDOM}};
  lineBuffer_4782 = _RAND_4789[7:0];
  _RAND_4790 = {1{`RANDOM}};
  lineBuffer_4783 = _RAND_4790[7:0];
  _RAND_4791 = {1{`RANDOM}};
  lineBuffer_4784 = _RAND_4791[7:0];
  _RAND_4792 = {1{`RANDOM}};
  lineBuffer_4785 = _RAND_4792[7:0];
  _RAND_4793 = {1{`RANDOM}};
  lineBuffer_4786 = _RAND_4793[7:0];
  _RAND_4794 = {1{`RANDOM}};
  lineBuffer_4787 = _RAND_4794[7:0];
  _RAND_4795 = {1{`RANDOM}};
  lineBuffer_4788 = _RAND_4795[7:0];
  _RAND_4796 = {1{`RANDOM}};
  lineBuffer_4789 = _RAND_4796[7:0];
  _RAND_4797 = {1{`RANDOM}};
  lineBuffer_4790 = _RAND_4797[7:0];
  _RAND_4798 = {1{`RANDOM}};
  lineBuffer_4791 = _RAND_4798[7:0];
  _RAND_4799 = {1{`RANDOM}};
  lineBuffer_4792 = _RAND_4799[7:0];
  _RAND_4800 = {1{`RANDOM}};
  lineBuffer_4793 = _RAND_4800[7:0];
  _RAND_4801 = {1{`RANDOM}};
  lineBuffer_4794 = _RAND_4801[7:0];
  _RAND_4802 = {1{`RANDOM}};
  lineBuffer_4795 = _RAND_4802[7:0];
  _RAND_4803 = {1{`RANDOM}};
  lineBuffer_4796 = _RAND_4803[7:0];
  _RAND_4804 = {1{`RANDOM}};
  lineBuffer_4797 = _RAND_4804[7:0];
  _RAND_4805 = {1{`RANDOM}};
  lineBuffer_4798 = _RAND_4805[7:0];
  _RAND_4806 = {1{`RANDOM}};
  lineBuffer_4799 = _RAND_4806[7:0];
  _RAND_4807 = {1{`RANDOM}};
  lineBuffer_4800 = _RAND_4807[7:0];
  _RAND_4808 = {1{`RANDOM}};
  lineBuffer_4801 = _RAND_4808[7:0];
  _RAND_4809 = {1{`RANDOM}};
  lineBuffer_4802 = _RAND_4809[7:0];
  _RAND_4810 = {1{`RANDOM}};
  lineBuffer_4803 = _RAND_4810[7:0];
  _RAND_4811 = {1{`RANDOM}};
  lineBuffer_4804 = _RAND_4811[7:0];
  _RAND_4812 = {1{`RANDOM}};
  lineBuffer_4805 = _RAND_4812[7:0];
  _RAND_4813 = {1{`RANDOM}};
  lineBuffer_4806 = _RAND_4813[7:0];
  _RAND_4814 = {1{`RANDOM}};
  lineBuffer_4807 = _RAND_4814[7:0];
  _RAND_4815 = {1{`RANDOM}};
  lineBuffer_4808 = _RAND_4815[7:0];
  _RAND_4816 = {1{`RANDOM}};
  lineBuffer_4809 = _RAND_4816[7:0];
  _RAND_4817 = {1{`RANDOM}};
  lineBuffer_4810 = _RAND_4817[7:0];
  _RAND_4818 = {1{`RANDOM}};
  lineBuffer_4811 = _RAND_4818[7:0];
  _RAND_4819 = {1{`RANDOM}};
  lineBuffer_4812 = _RAND_4819[7:0];
  _RAND_4820 = {1{`RANDOM}};
  lineBuffer_4813 = _RAND_4820[7:0];
  _RAND_4821 = {1{`RANDOM}};
  lineBuffer_4814 = _RAND_4821[7:0];
  _RAND_4822 = {1{`RANDOM}};
  lineBuffer_4815 = _RAND_4822[7:0];
  _RAND_4823 = {1{`RANDOM}};
  lineBuffer_4816 = _RAND_4823[7:0];
  _RAND_4824 = {1{`RANDOM}};
  lineBuffer_4817 = _RAND_4824[7:0];
  _RAND_4825 = {1{`RANDOM}};
  lineBuffer_4818 = _RAND_4825[7:0];
  _RAND_4826 = {1{`RANDOM}};
  lineBuffer_4819 = _RAND_4826[7:0];
  _RAND_4827 = {1{`RANDOM}};
  lineBuffer_4820 = _RAND_4827[7:0];
  _RAND_4828 = {1{`RANDOM}};
  lineBuffer_4821 = _RAND_4828[7:0];
  _RAND_4829 = {1{`RANDOM}};
  lineBuffer_4822 = _RAND_4829[7:0];
  _RAND_4830 = {1{`RANDOM}};
  lineBuffer_4823 = _RAND_4830[7:0];
  _RAND_4831 = {1{`RANDOM}};
  lineBuffer_4824 = _RAND_4831[7:0];
  _RAND_4832 = {1{`RANDOM}};
  lineBuffer_4825 = _RAND_4832[7:0];
  _RAND_4833 = {1{`RANDOM}};
  lineBuffer_4826 = _RAND_4833[7:0];
  _RAND_4834 = {1{`RANDOM}};
  lineBuffer_4827 = _RAND_4834[7:0];
  _RAND_4835 = {1{`RANDOM}};
  lineBuffer_4828 = _RAND_4835[7:0];
  _RAND_4836 = {1{`RANDOM}};
  lineBuffer_4829 = _RAND_4836[7:0];
  _RAND_4837 = {1{`RANDOM}};
  lineBuffer_4830 = _RAND_4837[7:0];
  _RAND_4838 = {1{`RANDOM}};
  lineBuffer_4831 = _RAND_4838[7:0];
  _RAND_4839 = {1{`RANDOM}};
  lineBuffer_4832 = _RAND_4839[7:0];
  _RAND_4840 = {1{`RANDOM}};
  lineBuffer_4833 = _RAND_4840[7:0];
  _RAND_4841 = {1{`RANDOM}};
  lineBuffer_4834 = _RAND_4841[7:0];
  _RAND_4842 = {1{`RANDOM}};
  lineBuffer_4835 = _RAND_4842[7:0];
  _RAND_4843 = {1{`RANDOM}};
  lineBuffer_4836 = _RAND_4843[7:0];
  _RAND_4844 = {1{`RANDOM}};
  lineBuffer_4837 = _RAND_4844[7:0];
  _RAND_4845 = {1{`RANDOM}};
  lineBuffer_4838 = _RAND_4845[7:0];
  _RAND_4846 = {1{`RANDOM}};
  lineBuffer_4839 = _RAND_4846[7:0];
  _RAND_4847 = {1{`RANDOM}};
  lineBuffer_4840 = _RAND_4847[7:0];
  _RAND_4848 = {1{`RANDOM}};
  lineBuffer_4841 = _RAND_4848[7:0];
  _RAND_4849 = {1{`RANDOM}};
  lineBuffer_4842 = _RAND_4849[7:0];
  _RAND_4850 = {1{`RANDOM}};
  lineBuffer_4843 = _RAND_4850[7:0];
  _RAND_4851 = {1{`RANDOM}};
  lineBuffer_4844 = _RAND_4851[7:0];
  _RAND_4852 = {1{`RANDOM}};
  lineBuffer_4845 = _RAND_4852[7:0];
  _RAND_4853 = {1{`RANDOM}};
  lineBuffer_4846 = _RAND_4853[7:0];
  _RAND_4854 = {1{`RANDOM}};
  lineBuffer_4847 = _RAND_4854[7:0];
  _RAND_4855 = {1{`RANDOM}};
  lineBuffer_4848 = _RAND_4855[7:0];
  _RAND_4856 = {1{`RANDOM}};
  lineBuffer_4849 = _RAND_4856[7:0];
  _RAND_4857 = {1{`RANDOM}};
  lineBuffer_4850 = _RAND_4857[7:0];
  _RAND_4858 = {1{`RANDOM}};
  lineBuffer_4851 = _RAND_4858[7:0];
  _RAND_4859 = {1{`RANDOM}};
  lineBuffer_4852 = _RAND_4859[7:0];
  _RAND_4860 = {1{`RANDOM}};
  lineBuffer_4853 = _RAND_4860[7:0];
  _RAND_4861 = {1{`RANDOM}};
  lineBuffer_4854 = _RAND_4861[7:0];
  _RAND_4862 = {1{`RANDOM}};
  lineBuffer_4855 = _RAND_4862[7:0];
  _RAND_4863 = {1{`RANDOM}};
  lineBuffer_4856 = _RAND_4863[7:0];
  _RAND_4864 = {1{`RANDOM}};
  lineBuffer_4857 = _RAND_4864[7:0];
  _RAND_4865 = {1{`RANDOM}};
  lineBuffer_4858 = _RAND_4865[7:0];
  _RAND_4866 = {1{`RANDOM}};
  lineBuffer_4859 = _RAND_4866[7:0];
  _RAND_4867 = {1{`RANDOM}};
  lineBuffer_4860 = _RAND_4867[7:0];
  _RAND_4868 = {1{`RANDOM}};
  lineBuffer_4861 = _RAND_4868[7:0];
  _RAND_4869 = {1{`RANDOM}};
  lineBuffer_4862 = _RAND_4869[7:0];
  _RAND_4870 = {1{`RANDOM}};
  lineBuffer_4863 = _RAND_4870[7:0];
  _RAND_4871 = {1{`RANDOM}};
  lineBuffer_4864 = _RAND_4871[7:0];
  _RAND_4872 = {1{`RANDOM}};
  lineBuffer_4865 = _RAND_4872[7:0];
  _RAND_4873 = {1{`RANDOM}};
  lineBuffer_4866 = _RAND_4873[7:0];
  _RAND_4874 = {1{`RANDOM}};
  lineBuffer_4867 = _RAND_4874[7:0];
  _RAND_4875 = {1{`RANDOM}};
  lineBuffer_4868 = _RAND_4875[7:0];
  _RAND_4876 = {1{`RANDOM}};
  lineBuffer_4869 = _RAND_4876[7:0];
  _RAND_4877 = {1{`RANDOM}};
  lineBuffer_4870 = _RAND_4877[7:0];
  _RAND_4878 = {1{`RANDOM}};
  lineBuffer_4871 = _RAND_4878[7:0];
  _RAND_4879 = {1{`RANDOM}};
  lineBuffer_4872 = _RAND_4879[7:0];
  _RAND_4880 = {1{`RANDOM}};
  lineBuffer_4873 = _RAND_4880[7:0];
  _RAND_4881 = {1{`RANDOM}};
  lineBuffer_4874 = _RAND_4881[7:0];
  _RAND_4882 = {1{`RANDOM}};
  lineBuffer_4875 = _RAND_4882[7:0];
  _RAND_4883 = {1{`RANDOM}};
  lineBuffer_4876 = _RAND_4883[7:0];
  _RAND_4884 = {1{`RANDOM}};
  lineBuffer_4877 = _RAND_4884[7:0];
  _RAND_4885 = {1{`RANDOM}};
  lineBuffer_4878 = _RAND_4885[7:0];
  _RAND_4886 = {1{`RANDOM}};
  lineBuffer_4879 = _RAND_4886[7:0];
  _RAND_4887 = {1{`RANDOM}};
  lineBuffer_4880 = _RAND_4887[7:0];
  _RAND_4888 = {1{`RANDOM}};
  lineBuffer_4881 = _RAND_4888[7:0];
  _RAND_4889 = {1{`RANDOM}};
  lineBuffer_4882 = _RAND_4889[7:0];
  _RAND_4890 = {1{`RANDOM}};
  lineBuffer_4883 = _RAND_4890[7:0];
  _RAND_4891 = {1{`RANDOM}};
  lineBuffer_4884 = _RAND_4891[7:0];
  _RAND_4892 = {1{`RANDOM}};
  lineBuffer_4885 = _RAND_4892[7:0];
  _RAND_4893 = {1{`RANDOM}};
  lineBuffer_4886 = _RAND_4893[7:0];
  _RAND_4894 = {1{`RANDOM}};
  lineBuffer_4887 = _RAND_4894[7:0];
  _RAND_4895 = {1{`RANDOM}};
  lineBuffer_4888 = _RAND_4895[7:0];
  _RAND_4896 = {1{`RANDOM}};
  lineBuffer_4889 = _RAND_4896[7:0];
  _RAND_4897 = {1{`RANDOM}};
  lineBuffer_4890 = _RAND_4897[7:0];
  _RAND_4898 = {1{`RANDOM}};
  lineBuffer_4891 = _RAND_4898[7:0];
  _RAND_4899 = {1{`RANDOM}};
  lineBuffer_4892 = _RAND_4899[7:0];
  _RAND_4900 = {1{`RANDOM}};
  lineBuffer_4893 = _RAND_4900[7:0];
  _RAND_4901 = {1{`RANDOM}};
  lineBuffer_4894 = _RAND_4901[7:0];
  _RAND_4902 = {1{`RANDOM}};
  lineBuffer_4895 = _RAND_4902[7:0];
  _RAND_4903 = {1{`RANDOM}};
  lineBuffer_4896 = _RAND_4903[7:0];
  _RAND_4904 = {1{`RANDOM}};
  lineBuffer_4897 = _RAND_4904[7:0];
  _RAND_4905 = {1{`RANDOM}};
  lineBuffer_4898 = _RAND_4905[7:0];
  _RAND_4906 = {1{`RANDOM}};
  lineBuffer_4899 = _RAND_4906[7:0];
  _RAND_4907 = {1{`RANDOM}};
  lineBuffer_4900 = _RAND_4907[7:0];
  _RAND_4908 = {1{`RANDOM}};
  lineBuffer_4901 = _RAND_4908[7:0];
  _RAND_4909 = {1{`RANDOM}};
  lineBuffer_4902 = _RAND_4909[7:0];
  _RAND_4910 = {1{`RANDOM}};
  lineBuffer_4903 = _RAND_4910[7:0];
  _RAND_4911 = {1{`RANDOM}};
  lineBuffer_4904 = _RAND_4911[7:0];
  _RAND_4912 = {1{`RANDOM}};
  lineBuffer_4905 = _RAND_4912[7:0];
  _RAND_4913 = {1{`RANDOM}};
  lineBuffer_4906 = _RAND_4913[7:0];
  _RAND_4914 = {1{`RANDOM}};
  lineBuffer_4907 = _RAND_4914[7:0];
  _RAND_4915 = {1{`RANDOM}};
  lineBuffer_4908 = _RAND_4915[7:0];
  _RAND_4916 = {1{`RANDOM}};
  lineBuffer_4909 = _RAND_4916[7:0];
  _RAND_4917 = {1{`RANDOM}};
  lineBuffer_4910 = _RAND_4917[7:0];
  _RAND_4918 = {1{`RANDOM}};
  lineBuffer_4911 = _RAND_4918[7:0];
  _RAND_4919 = {1{`RANDOM}};
  lineBuffer_4912 = _RAND_4919[7:0];
  _RAND_4920 = {1{`RANDOM}};
  lineBuffer_4913 = _RAND_4920[7:0];
  _RAND_4921 = {1{`RANDOM}};
  lineBuffer_4914 = _RAND_4921[7:0];
  _RAND_4922 = {1{`RANDOM}};
  lineBuffer_4915 = _RAND_4922[7:0];
  _RAND_4923 = {1{`RANDOM}};
  lineBuffer_4916 = _RAND_4923[7:0];
  _RAND_4924 = {1{`RANDOM}};
  lineBuffer_4917 = _RAND_4924[7:0];
  _RAND_4925 = {1{`RANDOM}};
  lineBuffer_4918 = _RAND_4925[7:0];
  _RAND_4926 = {1{`RANDOM}};
  lineBuffer_4919 = _RAND_4926[7:0];
  _RAND_4927 = {1{`RANDOM}};
  lineBuffer_4920 = _RAND_4927[7:0];
  _RAND_4928 = {1{`RANDOM}};
  lineBuffer_4921 = _RAND_4928[7:0];
  _RAND_4929 = {1{`RANDOM}};
  lineBuffer_4922 = _RAND_4929[7:0];
  _RAND_4930 = {1{`RANDOM}};
  lineBuffer_4923 = _RAND_4930[7:0];
  _RAND_4931 = {1{`RANDOM}};
  lineBuffer_4924 = _RAND_4931[7:0];
  _RAND_4932 = {1{`RANDOM}};
  lineBuffer_4925 = _RAND_4932[7:0];
  _RAND_4933 = {1{`RANDOM}};
  lineBuffer_4926 = _RAND_4933[7:0];
  _RAND_4934 = {1{`RANDOM}};
  lineBuffer_4927 = _RAND_4934[7:0];
  _RAND_4935 = {1{`RANDOM}};
  lineBuffer_4928 = _RAND_4935[7:0];
  _RAND_4936 = {1{`RANDOM}};
  lineBuffer_4929 = _RAND_4936[7:0];
  _RAND_4937 = {1{`RANDOM}};
  lineBuffer_4930 = _RAND_4937[7:0];
  _RAND_4938 = {1{`RANDOM}};
  lineBuffer_4931 = _RAND_4938[7:0];
  _RAND_4939 = {1{`RANDOM}};
  lineBuffer_4932 = _RAND_4939[7:0];
  _RAND_4940 = {1{`RANDOM}};
  lineBuffer_4933 = _RAND_4940[7:0];
  _RAND_4941 = {1{`RANDOM}};
  lineBuffer_4934 = _RAND_4941[7:0];
  _RAND_4942 = {1{`RANDOM}};
  lineBuffer_4935 = _RAND_4942[7:0];
  _RAND_4943 = {1{`RANDOM}};
  lineBuffer_4936 = _RAND_4943[7:0];
  _RAND_4944 = {1{`RANDOM}};
  lineBuffer_4937 = _RAND_4944[7:0];
  _RAND_4945 = {1{`RANDOM}};
  lineBuffer_4938 = _RAND_4945[7:0];
  _RAND_4946 = {1{`RANDOM}};
  lineBuffer_4939 = _RAND_4946[7:0];
  _RAND_4947 = {1{`RANDOM}};
  lineBuffer_4940 = _RAND_4947[7:0];
  _RAND_4948 = {1{`RANDOM}};
  lineBuffer_4941 = _RAND_4948[7:0];
  _RAND_4949 = {1{`RANDOM}};
  lineBuffer_4942 = _RAND_4949[7:0];
  _RAND_4950 = {1{`RANDOM}};
  lineBuffer_4943 = _RAND_4950[7:0];
  _RAND_4951 = {1{`RANDOM}};
  lineBuffer_4944 = _RAND_4951[7:0];
  _RAND_4952 = {1{`RANDOM}};
  lineBuffer_4945 = _RAND_4952[7:0];
  _RAND_4953 = {1{`RANDOM}};
  lineBuffer_4946 = _RAND_4953[7:0];
  _RAND_4954 = {1{`RANDOM}};
  lineBuffer_4947 = _RAND_4954[7:0];
  _RAND_4955 = {1{`RANDOM}};
  lineBuffer_4948 = _RAND_4955[7:0];
  _RAND_4956 = {1{`RANDOM}};
  lineBuffer_4949 = _RAND_4956[7:0];
  _RAND_4957 = {1{`RANDOM}};
  lineBuffer_4950 = _RAND_4957[7:0];
  _RAND_4958 = {1{`RANDOM}};
  lineBuffer_4951 = _RAND_4958[7:0];
  _RAND_4959 = {1{`RANDOM}};
  lineBuffer_4952 = _RAND_4959[7:0];
  _RAND_4960 = {1{`RANDOM}};
  lineBuffer_4953 = _RAND_4960[7:0];
  _RAND_4961 = {1{`RANDOM}};
  lineBuffer_4954 = _RAND_4961[7:0];
  _RAND_4962 = {1{`RANDOM}};
  lineBuffer_4955 = _RAND_4962[7:0];
  _RAND_4963 = {1{`RANDOM}};
  lineBuffer_4956 = _RAND_4963[7:0];
  _RAND_4964 = {1{`RANDOM}};
  lineBuffer_4957 = _RAND_4964[7:0];
  _RAND_4965 = {1{`RANDOM}};
  lineBuffer_4958 = _RAND_4965[7:0];
  _RAND_4966 = {1{`RANDOM}};
  lineBuffer_4959 = _RAND_4966[7:0];
  _RAND_4967 = {1{`RANDOM}};
  lineBuffer_4960 = _RAND_4967[7:0];
  _RAND_4968 = {1{`RANDOM}};
  lineBuffer_4961 = _RAND_4968[7:0];
  _RAND_4969 = {1{`RANDOM}};
  lineBuffer_4962 = _RAND_4969[7:0];
  _RAND_4970 = {1{`RANDOM}};
  lineBuffer_4963 = _RAND_4970[7:0];
  _RAND_4971 = {1{`RANDOM}};
  lineBuffer_4964 = _RAND_4971[7:0];
  _RAND_4972 = {1{`RANDOM}};
  lineBuffer_4965 = _RAND_4972[7:0];
  _RAND_4973 = {1{`RANDOM}};
  lineBuffer_4966 = _RAND_4973[7:0];
  _RAND_4974 = {1{`RANDOM}};
  lineBuffer_4967 = _RAND_4974[7:0];
  _RAND_4975 = {1{`RANDOM}};
  lineBuffer_4968 = _RAND_4975[7:0];
  _RAND_4976 = {1{`RANDOM}};
  lineBuffer_4969 = _RAND_4976[7:0];
  _RAND_4977 = {1{`RANDOM}};
  lineBuffer_4970 = _RAND_4977[7:0];
  _RAND_4978 = {1{`RANDOM}};
  lineBuffer_4971 = _RAND_4978[7:0];
  _RAND_4979 = {1{`RANDOM}};
  lineBuffer_4972 = _RAND_4979[7:0];
  _RAND_4980 = {1{`RANDOM}};
  lineBuffer_4973 = _RAND_4980[7:0];
  _RAND_4981 = {1{`RANDOM}};
  lineBuffer_4974 = _RAND_4981[7:0];
  _RAND_4982 = {1{`RANDOM}};
  lineBuffer_4975 = _RAND_4982[7:0];
  _RAND_4983 = {1{`RANDOM}};
  lineBuffer_4976 = _RAND_4983[7:0];
  _RAND_4984 = {1{`RANDOM}};
  lineBuffer_4977 = _RAND_4984[7:0];
  _RAND_4985 = {1{`RANDOM}};
  lineBuffer_4978 = _RAND_4985[7:0];
  _RAND_4986 = {1{`RANDOM}};
  lineBuffer_4979 = _RAND_4986[7:0];
  _RAND_4987 = {1{`RANDOM}};
  lineBuffer_4980 = _RAND_4987[7:0];
  _RAND_4988 = {1{`RANDOM}};
  lineBuffer_4981 = _RAND_4988[7:0];
  _RAND_4989 = {1{`RANDOM}};
  lineBuffer_4982 = _RAND_4989[7:0];
  _RAND_4990 = {1{`RANDOM}};
  lineBuffer_4983 = _RAND_4990[7:0];
  _RAND_4991 = {1{`RANDOM}};
  lineBuffer_4984 = _RAND_4991[7:0];
  _RAND_4992 = {1{`RANDOM}};
  lineBuffer_4985 = _RAND_4992[7:0];
  _RAND_4993 = {1{`RANDOM}};
  lineBuffer_4986 = _RAND_4993[7:0];
  _RAND_4994 = {1{`RANDOM}};
  lineBuffer_4987 = _RAND_4994[7:0];
  _RAND_4995 = {1{`RANDOM}};
  lineBuffer_4988 = _RAND_4995[7:0];
  _RAND_4996 = {1{`RANDOM}};
  lineBuffer_4989 = _RAND_4996[7:0];
  _RAND_4997 = {1{`RANDOM}};
  lineBuffer_4990 = _RAND_4997[7:0];
  _RAND_4998 = {1{`RANDOM}};
  lineBuffer_4991 = _RAND_4998[7:0];
  _RAND_4999 = {1{`RANDOM}};
  lineBuffer_4992 = _RAND_4999[7:0];
  _RAND_5000 = {1{`RANDOM}};
  lineBuffer_4993 = _RAND_5000[7:0];
  _RAND_5001 = {1{`RANDOM}};
  lineBuffer_4994 = _RAND_5001[7:0];
  _RAND_5002 = {1{`RANDOM}};
  lineBuffer_4995 = _RAND_5002[7:0];
  _RAND_5003 = {1{`RANDOM}};
  lineBuffer_4996 = _RAND_5003[7:0];
  _RAND_5004 = {1{`RANDOM}};
  lineBuffer_4997 = _RAND_5004[7:0];
  _RAND_5005 = {1{`RANDOM}};
  lineBuffer_4998 = _RAND_5005[7:0];
  _RAND_5006 = {1{`RANDOM}};
  lineBuffer_4999 = _RAND_5006[7:0];
  _RAND_5007 = {1{`RANDOM}};
  lineBuffer_5000 = _RAND_5007[7:0];
  _RAND_5008 = {1{`RANDOM}};
  lineBuffer_5001 = _RAND_5008[7:0];
  _RAND_5009 = {1{`RANDOM}};
  lineBuffer_5002 = _RAND_5009[7:0];
  _RAND_5010 = {1{`RANDOM}};
  lineBuffer_5003 = _RAND_5010[7:0];
  _RAND_5011 = {1{`RANDOM}};
  lineBuffer_5004 = _RAND_5011[7:0];
  _RAND_5012 = {1{`RANDOM}};
  lineBuffer_5005 = _RAND_5012[7:0];
  _RAND_5013 = {1{`RANDOM}};
  lineBuffer_5006 = _RAND_5013[7:0];
  _RAND_5014 = {1{`RANDOM}};
  lineBuffer_5007 = _RAND_5014[7:0];
  _RAND_5015 = {1{`RANDOM}};
  lineBuffer_5008 = _RAND_5015[7:0];
  _RAND_5016 = {1{`RANDOM}};
  lineBuffer_5009 = _RAND_5016[7:0];
  _RAND_5017 = {1{`RANDOM}};
  lineBuffer_5010 = _RAND_5017[7:0];
  _RAND_5018 = {1{`RANDOM}};
  lineBuffer_5011 = _RAND_5018[7:0];
  _RAND_5019 = {1{`RANDOM}};
  lineBuffer_5012 = _RAND_5019[7:0];
  _RAND_5020 = {1{`RANDOM}};
  lineBuffer_5013 = _RAND_5020[7:0];
  _RAND_5021 = {1{`RANDOM}};
  lineBuffer_5014 = _RAND_5021[7:0];
  _RAND_5022 = {1{`RANDOM}};
  lineBuffer_5015 = _RAND_5022[7:0];
  _RAND_5023 = {1{`RANDOM}};
  lineBuffer_5016 = _RAND_5023[7:0];
  _RAND_5024 = {1{`RANDOM}};
  lineBuffer_5017 = _RAND_5024[7:0];
  _RAND_5025 = {1{`RANDOM}};
  lineBuffer_5018 = _RAND_5025[7:0];
  _RAND_5026 = {1{`RANDOM}};
  lineBuffer_5019 = _RAND_5026[7:0];
  _RAND_5027 = {1{`RANDOM}};
  lineBuffer_5020 = _RAND_5027[7:0];
  _RAND_5028 = {1{`RANDOM}};
  lineBuffer_5021 = _RAND_5028[7:0];
  _RAND_5029 = {1{`RANDOM}};
  lineBuffer_5022 = _RAND_5029[7:0];
  _RAND_5030 = {1{`RANDOM}};
  lineBuffer_5023 = _RAND_5030[7:0];
  _RAND_5031 = {1{`RANDOM}};
  lineBuffer_5024 = _RAND_5031[7:0];
  _RAND_5032 = {1{`RANDOM}};
  lineBuffer_5025 = _RAND_5032[7:0];
  _RAND_5033 = {1{`RANDOM}};
  lineBuffer_5026 = _RAND_5033[7:0];
  _RAND_5034 = {1{`RANDOM}};
  lineBuffer_5027 = _RAND_5034[7:0];
  _RAND_5035 = {1{`RANDOM}};
  lineBuffer_5028 = _RAND_5035[7:0];
  _RAND_5036 = {1{`RANDOM}};
  lineBuffer_5029 = _RAND_5036[7:0];
  _RAND_5037 = {1{`RANDOM}};
  lineBuffer_5030 = _RAND_5037[7:0];
  _RAND_5038 = {1{`RANDOM}};
  lineBuffer_5031 = _RAND_5038[7:0];
  _RAND_5039 = {1{`RANDOM}};
  lineBuffer_5032 = _RAND_5039[7:0];
  _RAND_5040 = {1{`RANDOM}};
  lineBuffer_5033 = _RAND_5040[7:0];
  _RAND_5041 = {1{`RANDOM}};
  lineBuffer_5034 = _RAND_5041[7:0];
  _RAND_5042 = {1{`RANDOM}};
  lineBuffer_5035 = _RAND_5042[7:0];
  _RAND_5043 = {1{`RANDOM}};
  lineBuffer_5036 = _RAND_5043[7:0];
  _RAND_5044 = {1{`RANDOM}};
  lineBuffer_5037 = _RAND_5044[7:0];
  _RAND_5045 = {1{`RANDOM}};
  lineBuffer_5038 = _RAND_5045[7:0];
  _RAND_5046 = {1{`RANDOM}};
  lineBuffer_5039 = _RAND_5046[7:0];
  _RAND_5047 = {1{`RANDOM}};
  lineBuffer_5040 = _RAND_5047[7:0];
  _RAND_5048 = {1{`RANDOM}};
  lineBuffer_5041 = _RAND_5048[7:0];
  _RAND_5049 = {1{`RANDOM}};
  lineBuffer_5042 = _RAND_5049[7:0];
  _RAND_5050 = {1{`RANDOM}};
  lineBuffer_5043 = _RAND_5050[7:0];
  _RAND_5051 = {1{`RANDOM}};
  lineBuffer_5044 = _RAND_5051[7:0];
  _RAND_5052 = {1{`RANDOM}};
  lineBuffer_5045 = _RAND_5052[7:0];
  _RAND_5053 = {1{`RANDOM}};
  lineBuffer_5046 = _RAND_5053[7:0];
  _RAND_5054 = {1{`RANDOM}};
  lineBuffer_5047 = _RAND_5054[7:0];
  _RAND_5055 = {1{`RANDOM}};
  lineBuffer_5048 = _RAND_5055[7:0];
  _RAND_5056 = {1{`RANDOM}};
  lineBuffer_5049 = _RAND_5056[7:0];
  _RAND_5057 = {1{`RANDOM}};
  lineBuffer_5050 = _RAND_5057[7:0];
  _RAND_5058 = {1{`RANDOM}};
  lineBuffer_5051 = _RAND_5058[7:0];
  _RAND_5059 = {1{`RANDOM}};
  lineBuffer_5052 = _RAND_5059[7:0];
  _RAND_5060 = {1{`RANDOM}};
  lineBuffer_5053 = _RAND_5060[7:0];
  _RAND_5061 = {1{`RANDOM}};
  lineBuffer_5054 = _RAND_5061[7:0];
  _RAND_5062 = {1{`RANDOM}};
  lineBuffer_5055 = _RAND_5062[7:0];
  _RAND_5063 = {1{`RANDOM}};
  lineBuffer_5056 = _RAND_5063[7:0];
  _RAND_5064 = {1{`RANDOM}};
  lineBuffer_5057 = _RAND_5064[7:0];
  _RAND_5065 = {1{`RANDOM}};
  lineBuffer_5058 = _RAND_5065[7:0];
  _RAND_5066 = {1{`RANDOM}};
  lineBuffer_5059 = _RAND_5066[7:0];
  _RAND_5067 = {1{`RANDOM}};
  lineBuffer_5060 = _RAND_5067[7:0];
  _RAND_5068 = {1{`RANDOM}};
  lineBuffer_5061 = _RAND_5068[7:0];
  _RAND_5069 = {1{`RANDOM}};
  lineBuffer_5062 = _RAND_5069[7:0];
  _RAND_5070 = {1{`RANDOM}};
  lineBuffer_5063 = _RAND_5070[7:0];
  _RAND_5071 = {1{`RANDOM}};
  lineBuffer_5064 = _RAND_5071[7:0];
  _RAND_5072 = {1{`RANDOM}};
  lineBuffer_5065 = _RAND_5072[7:0];
  _RAND_5073 = {1{`RANDOM}};
  lineBuffer_5066 = _RAND_5073[7:0];
  _RAND_5074 = {1{`RANDOM}};
  lineBuffer_5067 = _RAND_5074[7:0];
  _RAND_5075 = {1{`RANDOM}};
  lineBuffer_5068 = _RAND_5075[7:0];
  _RAND_5076 = {1{`RANDOM}};
  lineBuffer_5069 = _RAND_5076[7:0];
  _RAND_5077 = {1{`RANDOM}};
  lineBuffer_5070 = _RAND_5077[7:0];
  _RAND_5078 = {1{`RANDOM}};
  lineBuffer_5071 = _RAND_5078[7:0];
  _RAND_5079 = {1{`RANDOM}};
  lineBuffer_5072 = _RAND_5079[7:0];
  _RAND_5080 = {1{`RANDOM}};
  lineBuffer_5073 = _RAND_5080[7:0];
  _RAND_5081 = {1{`RANDOM}};
  lineBuffer_5074 = _RAND_5081[7:0];
  _RAND_5082 = {1{`RANDOM}};
  lineBuffer_5075 = _RAND_5082[7:0];
  _RAND_5083 = {1{`RANDOM}};
  lineBuffer_5076 = _RAND_5083[7:0];
  _RAND_5084 = {1{`RANDOM}};
  lineBuffer_5077 = _RAND_5084[7:0];
  _RAND_5085 = {1{`RANDOM}};
  lineBuffer_5078 = _RAND_5085[7:0];
  _RAND_5086 = {1{`RANDOM}};
  lineBuffer_5079 = _RAND_5086[7:0];
  _RAND_5087 = {1{`RANDOM}};
  lineBuffer_5080 = _RAND_5087[7:0];
  _RAND_5088 = {1{`RANDOM}};
  lineBuffer_5081 = _RAND_5088[7:0];
  _RAND_5089 = {1{`RANDOM}};
  lineBuffer_5082 = _RAND_5089[7:0];
  _RAND_5090 = {1{`RANDOM}};
  lineBuffer_5083 = _RAND_5090[7:0];
  _RAND_5091 = {1{`RANDOM}};
  lineBuffer_5084 = _RAND_5091[7:0];
  _RAND_5092 = {1{`RANDOM}};
  lineBuffer_5085 = _RAND_5092[7:0];
  _RAND_5093 = {1{`RANDOM}};
  lineBuffer_5086 = _RAND_5093[7:0];
  _RAND_5094 = {1{`RANDOM}};
  lineBuffer_5087 = _RAND_5094[7:0];
  _RAND_5095 = {1{`RANDOM}};
  lineBuffer_5088 = _RAND_5095[7:0];
  _RAND_5096 = {1{`RANDOM}};
  lineBuffer_5089 = _RAND_5096[7:0];
  _RAND_5097 = {1{`RANDOM}};
  lineBuffer_5090 = _RAND_5097[7:0];
  _RAND_5098 = {1{`RANDOM}};
  lineBuffer_5091 = _RAND_5098[7:0];
  _RAND_5099 = {1{`RANDOM}};
  lineBuffer_5092 = _RAND_5099[7:0];
  _RAND_5100 = {1{`RANDOM}};
  lineBuffer_5093 = _RAND_5100[7:0];
  _RAND_5101 = {1{`RANDOM}};
  lineBuffer_5094 = _RAND_5101[7:0];
  _RAND_5102 = {1{`RANDOM}};
  lineBuffer_5095 = _RAND_5102[7:0];
  _RAND_5103 = {1{`RANDOM}};
  lineBuffer_5096 = _RAND_5103[7:0];
  _RAND_5104 = {1{`RANDOM}};
  lineBuffer_5097 = _RAND_5104[7:0];
  _RAND_5105 = {1{`RANDOM}};
  lineBuffer_5098 = _RAND_5105[7:0];
  _RAND_5106 = {1{`RANDOM}};
  lineBuffer_5099 = _RAND_5106[7:0];
  _RAND_5107 = {1{`RANDOM}};
  lineBuffer_5100 = _RAND_5107[7:0];
  _RAND_5108 = {1{`RANDOM}};
  lineBuffer_5101 = _RAND_5108[7:0];
  _RAND_5109 = {1{`RANDOM}};
  lineBuffer_5102 = _RAND_5109[7:0];
  _RAND_5110 = {1{`RANDOM}};
  lineBuffer_5103 = _RAND_5110[7:0];
  _RAND_5111 = {1{`RANDOM}};
  lineBuffer_5104 = _RAND_5111[7:0];
  _RAND_5112 = {1{`RANDOM}};
  lineBuffer_5105 = _RAND_5112[7:0];
  _RAND_5113 = {1{`RANDOM}};
  lineBuffer_5106 = _RAND_5113[7:0];
  _RAND_5114 = {1{`RANDOM}};
  lineBuffer_5107 = _RAND_5114[7:0];
  _RAND_5115 = {1{`RANDOM}};
  lineBuffer_5108 = _RAND_5115[7:0];
  _RAND_5116 = {1{`RANDOM}};
  lineBuffer_5109 = _RAND_5116[7:0];
  _RAND_5117 = {1{`RANDOM}};
  lineBuffer_5110 = _RAND_5117[7:0];
  _RAND_5118 = {1{`RANDOM}};
  lineBuffer_5111 = _RAND_5118[7:0];
  _RAND_5119 = {1{`RANDOM}};
  lineBuffer_5112 = _RAND_5119[7:0];
  _RAND_5120 = {1{`RANDOM}};
  lineBuffer_5113 = _RAND_5120[7:0];
  _RAND_5121 = {1{`RANDOM}};
  lineBuffer_5114 = _RAND_5121[7:0];
  _RAND_5122 = {1{`RANDOM}};
  lineBuffer_5115 = _RAND_5122[7:0];
  _RAND_5123 = {1{`RANDOM}};
  lineBuffer_5116 = _RAND_5123[7:0];
  _RAND_5124 = {1{`RANDOM}};
  lineBuffer_5117 = _RAND_5124[7:0];
  _RAND_5125 = {1{`RANDOM}};
  lineBuffer_5118 = _RAND_5125[7:0];
  _RAND_5126 = {1{`RANDOM}};
  lineBuffer_5119 = _RAND_5126[7:0];
  _RAND_5127 = {1{`RANDOM}};
  lineBuffer_5120 = _RAND_5127[7:0];
  _RAND_5128 = {1{`RANDOM}};
  lineBuffer_5121 = _RAND_5128[7:0];
  _RAND_5129 = {1{`RANDOM}};
  lineBuffer_5122 = _RAND_5129[7:0];
  _RAND_5130 = {1{`RANDOM}};
  lineBuffer_5123 = _RAND_5130[7:0];
  _RAND_5131 = {1{`RANDOM}};
  lineBuffer_5124 = _RAND_5131[7:0];
  _RAND_5132 = {1{`RANDOM}};
  lineBuffer_5125 = _RAND_5132[7:0];
  _RAND_5133 = {1{`RANDOM}};
  lineBuffer_5126 = _RAND_5133[7:0];
  _RAND_5134 = {1{`RANDOM}};
  lineBuffer_5127 = _RAND_5134[7:0];
  _RAND_5135 = {1{`RANDOM}};
  lineBuffer_5128 = _RAND_5135[7:0];
  _RAND_5136 = {1{`RANDOM}};
  lineBuffer_5129 = _RAND_5136[7:0];
  _RAND_5137 = {1{`RANDOM}};
  lineBuffer_5130 = _RAND_5137[7:0];
  _RAND_5138 = {1{`RANDOM}};
  lineBuffer_5131 = _RAND_5138[7:0];
  _RAND_5139 = {1{`RANDOM}};
  lineBuffer_5132 = _RAND_5139[7:0];
  _RAND_5140 = {1{`RANDOM}};
  lineBuffer_5133 = _RAND_5140[7:0];
  _RAND_5141 = {1{`RANDOM}};
  lineBuffer_5134 = _RAND_5141[7:0];
  _RAND_5142 = {1{`RANDOM}};
  lineBuffer_5135 = _RAND_5142[7:0];
  _RAND_5143 = {1{`RANDOM}};
  lineBuffer_5136 = _RAND_5143[7:0];
  _RAND_5144 = {1{`RANDOM}};
  lineBuffer_5137 = _RAND_5144[7:0];
  _RAND_5145 = {1{`RANDOM}};
  lineBuffer_5138 = _RAND_5145[7:0];
  _RAND_5146 = {1{`RANDOM}};
  lineBuffer_5139 = _RAND_5146[7:0];
  _RAND_5147 = {1{`RANDOM}};
  lineBuffer_5140 = _RAND_5147[7:0];
  _RAND_5148 = {1{`RANDOM}};
  lineBuffer_5141 = _RAND_5148[7:0];
  _RAND_5149 = {1{`RANDOM}};
  lineBuffer_5142 = _RAND_5149[7:0];
  _RAND_5150 = {1{`RANDOM}};
  lineBuffer_5143 = _RAND_5150[7:0];
  _RAND_5151 = {1{`RANDOM}};
  lineBuffer_5144 = _RAND_5151[7:0];
  _RAND_5152 = {1{`RANDOM}};
  lineBuffer_5145 = _RAND_5152[7:0];
  _RAND_5153 = {1{`RANDOM}};
  lineBuffer_5146 = _RAND_5153[7:0];
  _RAND_5154 = {1{`RANDOM}};
  lineBuffer_5147 = _RAND_5154[7:0];
  _RAND_5155 = {1{`RANDOM}};
  lineBuffer_5148 = _RAND_5155[7:0];
  _RAND_5156 = {1{`RANDOM}};
  lineBuffer_5149 = _RAND_5156[7:0];
  _RAND_5157 = {1{`RANDOM}};
  lineBuffer_5150 = _RAND_5157[7:0];
  _RAND_5158 = {1{`RANDOM}};
  lineBuffer_5151 = _RAND_5158[7:0];
  _RAND_5159 = {1{`RANDOM}};
  lineBuffer_5152 = _RAND_5159[7:0];
  _RAND_5160 = {1{`RANDOM}};
  lineBuffer_5153 = _RAND_5160[7:0];
  _RAND_5161 = {1{`RANDOM}};
  lineBuffer_5154 = _RAND_5161[7:0];
  _RAND_5162 = {1{`RANDOM}};
  lineBuffer_5155 = _RAND_5162[7:0];
  _RAND_5163 = {1{`RANDOM}};
  lineBuffer_5156 = _RAND_5163[7:0];
  _RAND_5164 = {1{`RANDOM}};
  lineBuffer_5157 = _RAND_5164[7:0];
  _RAND_5165 = {1{`RANDOM}};
  lineBuffer_5158 = _RAND_5165[7:0];
  _RAND_5166 = {1{`RANDOM}};
  lineBuffer_5159 = _RAND_5166[7:0];
  _RAND_5167 = {1{`RANDOM}};
  lineBuffer_5160 = _RAND_5167[7:0];
  _RAND_5168 = {1{`RANDOM}};
  lineBuffer_5161 = _RAND_5168[7:0];
  _RAND_5169 = {1{`RANDOM}};
  lineBuffer_5162 = _RAND_5169[7:0];
  _RAND_5170 = {1{`RANDOM}};
  lineBuffer_5163 = _RAND_5170[7:0];
  _RAND_5171 = {1{`RANDOM}};
  lineBuffer_5164 = _RAND_5171[7:0];
  _RAND_5172 = {1{`RANDOM}};
  lineBuffer_5165 = _RAND_5172[7:0];
  _RAND_5173 = {1{`RANDOM}};
  lineBuffer_5166 = _RAND_5173[7:0];
  _RAND_5174 = {1{`RANDOM}};
  lineBuffer_5167 = _RAND_5174[7:0];
  _RAND_5175 = {1{`RANDOM}};
  lineBuffer_5168 = _RAND_5175[7:0];
  _RAND_5176 = {1{`RANDOM}};
  lineBuffer_5169 = _RAND_5176[7:0];
  _RAND_5177 = {1{`RANDOM}};
  lineBuffer_5170 = _RAND_5177[7:0];
  _RAND_5178 = {1{`RANDOM}};
  lineBuffer_5171 = _RAND_5178[7:0];
  _RAND_5179 = {1{`RANDOM}};
  lineBuffer_5172 = _RAND_5179[7:0];
  _RAND_5180 = {1{`RANDOM}};
  lineBuffer_5173 = _RAND_5180[7:0];
  _RAND_5181 = {1{`RANDOM}};
  lineBuffer_5174 = _RAND_5181[7:0];
  _RAND_5182 = {1{`RANDOM}};
  lineBuffer_5175 = _RAND_5182[7:0];
  _RAND_5183 = {1{`RANDOM}};
  lineBuffer_5176 = _RAND_5183[7:0];
  _RAND_5184 = {1{`RANDOM}};
  lineBuffer_5177 = _RAND_5184[7:0];
  _RAND_5185 = {1{`RANDOM}};
  lineBuffer_5178 = _RAND_5185[7:0];
  _RAND_5186 = {1{`RANDOM}};
  lineBuffer_5179 = _RAND_5186[7:0];
  _RAND_5187 = {1{`RANDOM}};
  lineBuffer_5180 = _RAND_5187[7:0];
  _RAND_5188 = {1{`RANDOM}};
  lineBuffer_5181 = _RAND_5188[7:0];
  _RAND_5189 = {1{`RANDOM}};
  lineBuffer_5182 = _RAND_5189[7:0];
  _RAND_5190 = {1{`RANDOM}};
  lineBuffer_5183 = _RAND_5190[7:0];
  _RAND_5191 = {1{`RANDOM}};
  lineBuffer_5184 = _RAND_5191[7:0];
  _RAND_5192 = {1{`RANDOM}};
  lineBuffer_5185 = _RAND_5192[7:0];
  _RAND_5193 = {1{`RANDOM}};
  lineBuffer_5186 = _RAND_5193[7:0];
  _RAND_5194 = {1{`RANDOM}};
  lineBuffer_5187 = _RAND_5194[7:0];
  _RAND_5195 = {1{`RANDOM}};
  lineBuffer_5188 = _RAND_5195[7:0];
  _RAND_5196 = {1{`RANDOM}};
  lineBuffer_5189 = _RAND_5196[7:0];
  _RAND_5197 = {1{`RANDOM}};
  lineBuffer_5190 = _RAND_5197[7:0];
  _RAND_5198 = {1{`RANDOM}};
  lineBuffer_5191 = _RAND_5198[7:0];
  _RAND_5199 = {1{`RANDOM}};
  lineBuffer_5192 = _RAND_5199[7:0];
  _RAND_5200 = {1{`RANDOM}};
  lineBuffer_5193 = _RAND_5200[7:0];
  _RAND_5201 = {1{`RANDOM}};
  lineBuffer_5194 = _RAND_5201[7:0];
  _RAND_5202 = {1{`RANDOM}};
  lineBuffer_5195 = _RAND_5202[7:0];
  _RAND_5203 = {1{`RANDOM}};
  lineBuffer_5196 = _RAND_5203[7:0];
  _RAND_5204 = {1{`RANDOM}};
  lineBuffer_5197 = _RAND_5204[7:0];
  _RAND_5205 = {1{`RANDOM}};
  lineBuffer_5198 = _RAND_5205[7:0];
  _RAND_5206 = {1{`RANDOM}};
  lineBuffer_5199 = _RAND_5206[7:0];
  _RAND_5207 = {1{`RANDOM}};
  lineBuffer_5200 = _RAND_5207[7:0];
  _RAND_5208 = {1{`RANDOM}};
  lineBuffer_5201 = _RAND_5208[7:0];
  _RAND_5209 = {1{`RANDOM}};
  lineBuffer_5202 = _RAND_5209[7:0];
  _RAND_5210 = {1{`RANDOM}};
  lineBuffer_5203 = _RAND_5210[7:0];
  _RAND_5211 = {1{`RANDOM}};
  lineBuffer_5204 = _RAND_5211[7:0];
  _RAND_5212 = {1{`RANDOM}};
  lineBuffer_5205 = _RAND_5212[7:0];
  _RAND_5213 = {1{`RANDOM}};
  lineBuffer_5206 = _RAND_5213[7:0];
  _RAND_5214 = {1{`RANDOM}};
  lineBuffer_5207 = _RAND_5214[7:0];
  _RAND_5215 = {1{`RANDOM}};
  lineBuffer_5208 = _RAND_5215[7:0];
  _RAND_5216 = {1{`RANDOM}};
  lineBuffer_5209 = _RAND_5216[7:0];
  _RAND_5217 = {1{`RANDOM}};
  lineBuffer_5210 = _RAND_5217[7:0];
  _RAND_5218 = {1{`RANDOM}};
  lineBuffer_5211 = _RAND_5218[7:0];
  _RAND_5219 = {1{`RANDOM}};
  lineBuffer_5212 = _RAND_5219[7:0];
  _RAND_5220 = {1{`RANDOM}};
  lineBuffer_5213 = _RAND_5220[7:0];
  _RAND_5221 = {1{`RANDOM}};
  lineBuffer_5214 = _RAND_5221[7:0];
  _RAND_5222 = {1{`RANDOM}};
  lineBuffer_5215 = _RAND_5222[7:0];
  _RAND_5223 = {1{`RANDOM}};
  lineBuffer_5216 = _RAND_5223[7:0];
  _RAND_5224 = {1{`RANDOM}};
  lineBuffer_5217 = _RAND_5224[7:0];
  _RAND_5225 = {1{`RANDOM}};
  lineBuffer_5218 = _RAND_5225[7:0];
  _RAND_5226 = {1{`RANDOM}};
  lineBuffer_5219 = _RAND_5226[7:0];
  _RAND_5227 = {1{`RANDOM}};
  lineBuffer_5220 = _RAND_5227[7:0];
  _RAND_5228 = {1{`RANDOM}};
  lineBuffer_5221 = _RAND_5228[7:0];
  _RAND_5229 = {1{`RANDOM}};
  lineBuffer_5222 = _RAND_5229[7:0];
  _RAND_5230 = {1{`RANDOM}};
  lineBuffer_5223 = _RAND_5230[7:0];
  _RAND_5231 = {1{`RANDOM}};
  lineBuffer_5224 = _RAND_5231[7:0];
  _RAND_5232 = {1{`RANDOM}};
  lineBuffer_5225 = _RAND_5232[7:0];
  _RAND_5233 = {1{`RANDOM}};
  lineBuffer_5226 = _RAND_5233[7:0];
  _RAND_5234 = {1{`RANDOM}};
  lineBuffer_5227 = _RAND_5234[7:0];
  _RAND_5235 = {1{`RANDOM}};
  lineBuffer_5228 = _RAND_5235[7:0];
  _RAND_5236 = {1{`RANDOM}};
  lineBuffer_5229 = _RAND_5236[7:0];
  _RAND_5237 = {1{`RANDOM}};
  lineBuffer_5230 = _RAND_5237[7:0];
  _RAND_5238 = {1{`RANDOM}};
  lineBuffer_5231 = _RAND_5238[7:0];
  _RAND_5239 = {1{`RANDOM}};
  lineBuffer_5232 = _RAND_5239[7:0];
  _RAND_5240 = {1{`RANDOM}};
  lineBuffer_5233 = _RAND_5240[7:0];
  _RAND_5241 = {1{`RANDOM}};
  lineBuffer_5234 = _RAND_5241[7:0];
  _RAND_5242 = {1{`RANDOM}};
  lineBuffer_5235 = _RAND_5242[7:0];
  _RAND_5243 = {1{`RANDOM}};
  lineBuffer_5236 = _RAND_5243[7:0];
  _RAND_5244 = {1{`RANDOM}};
  lineBuffer_5237 = _RAND_5244[7:0];
  _RAND_5245 = {1{`RANDOM}};
  lineBuffer_5238 = _RAND_5245[7:0];
  _RAND_5246 = {1{`RANDOM}};
  lineBuffer_5239 = _RAND_5246[7:0];
  _RAND_5247 = {1{`RANDOM}};
  lineBuffer_5240 = _RAND_5247[7:0];
  _RAND_5248 = {1{`RANDOM}};
  lineBuffer_5241 = _RAND_5248[7:0];
  _RAND_5249 = {1{`RANDOM}};
  lineBuffer_5242 = _RAND_5249[7:0];
  _RAND_5250 = {1{`RANDOM}};
  lineBuffer_5243 = _RAND_5250[7:0];
  _RAND_5251 = {1{`RANDOM}};
  lineBuffer_5244 = _RAND_5251[7:0];
  _RAND_5252 = {1{`RANDOM}};
  lineBuffer_5245 = _RAND_5252[7:0];
  _RAND_5253 = {1{`RANDOM}};
  lineBuffer_5246 = _RAND_5253[7:0];
  _RAND_5254 = {1{`RANDOM}};
  lineBuffer_5247 = _RAND_5254[7:0];
  _RAND_5255 = {1{`RANDOM}};
  lineBuffer_5248 = _RAND_5255[7:0];
  _RAND_5256 = {1{`RANDOM}};
  lineBuffer_5249 = _RAND_5256[7:0];
  _RAND_5257 = {1{`RANDOM}};
  lineBuffer_5250 = _RAND_5257[7:0];
  _RAND_5258 = {1{`RANDOM}};
  lineBuffer_5251 = _RAND_5258[7:0];
  _RAND_5259 = {1{`RANDOM}};
  lineBuffer_5252 = _RAND_5259[7:0];
  _RAND_5260 = {1{`RANDOM}};
  lineBuffer_5253 = _RAND_5260[7:0];
  _RAND_5261 = {1{`RANDOM}};
  lineBuffer_5254 = _RAND_5261[7:0];
  _RAND_5262 = {1{`RANDOM}};
  lineBuffer_5255 = _RAND_5262[7:0];
  _RAND_5263 = {1{`RANDOM}};
  lineBuffer_5256 = _RAND_5263[7:0];
  _RAND_5264 = {1{`RANDOM}};
  lineBuffer_5257 = _RAND_5264[7:0];
  _RAND_5265 = {1{`RANDOM}};
  lineBuffer_5258 = _RAND_5265[7:0];
  _RAND_5266 = {1{`RANDOM}};
  lineBuffer_5259 = _RAND_5266[7:0];
  _RAND_5267 = {1{`RANDOM}};
  lineBuffer_5260 = _RAND_5267[7:0];
  _RAND_5268 = {1{`RANDOM}};
  lineBuffer_5261 = _RAND_5268[7:0];
  _RAND_5269 = {1{`RANDOM}};
  lineBuffer_5262 = _RAND_5269[7:0];
  _RAND_5270 = {1{`RANDOM}};
  lineBuffer_5263 = _RAND_5270[7:0];
  _RAND_5271 = {1{`RANDOM}};
  lineBuffer_5264 = _RAND_5271[7:0];
  _RAND_5272 = {1{`RANDOM}};
  lineBuffer_5265 = _RAND_5272[7:0];
  _RAND_5273 = {1{`RANDOM}};
  lineBuffer_5266 = _RAND_5273[7:0];
  _RAND_5274 = {1{`RANDOM}};
  lineBuffer_5267 = _RAND_5274[7:0];
  _RAND_5275 = {1{`RANDOM}};
  lineBuffer_5268 = _RAND_5275[7:0];
  _RAND_5276 = {1{`RANDOM}};
  lineBuffer_5269 = _RAND_5276[7:0];
  _RAND_5277 = {1{`RANDOM}};
  lineBuffer_5270 = _RAND_5277[7:0];
  _RAND_5278 = {1{`RANDOM}};
  lineBuffer_5271 = _RAND_5278[7:0];
  _RAND_5279 = {1{`RANDOM}};
  lineBuffer_5272 = _RAND_5279[7:0];
  _RAND_5280 = {1{`RANDOM}};
  lineBuffer_5273 = _RAND_5280[7:0];
  _RAND_5281 = {1{`RANDOM}};
  lineBuffer_5274 = _RAND_5281[7:0];
  _RAND_5282 = {1{`RANDOM}};
  lineBuffer_5275 = _RAND_5282[7:0];
  _RAND_5283 = {1{`RANDOM}};
  lineBuffer_5276 = _RAND_5283[7:0];
  _RAND_5284 = {1{`RANDOM}};
  lineBuffer_5277 = _RAND_5284[7:0];
  _RAND_5285 = {1{`RANDOM}};
  lineBuffer_5278 = _RAND_5285[7:0];
  _RAND_5286 = {1{`RANDOM}};
  lineBuffer_5279 = _RAND_5286[7:0];
  _RAND_5287 = {1{`RANDOM}};
  lineBuffer_5280 = _RAND_5287[7:0];
  _RAND_5288 = {1{`RANDOM}};
  lineBuffer_5281 = _RAND_5288[7:0];
  _RAND_5289 = {1{`RANDOM}};
  lineBuffer_5282 = _RAND_5289[7:0];
  _RAND_5290 = {1{`RANDOM}};
  lineBuffer_5283 = _RAND_5290[7:0];
  _RAND_5291 = {1{`RANDOM}};
  lineBuffer_5284 = _RAND_5291[7:0];
  _RAND_5292 = {1{`RANDOM}};
  lineBuffer_5285 = _RAND_5292[7:0];
  _RAND_5293 = {1{`RANDOM}};
  lineBuffer_5286 = _RAND_5293[7:0];
  _RAND_5294 = {1{`RANDOM}};
  lineBuffer_5287 = _RAND_5294[7:0];
  _RAND_5295 = {1{`RANDOM}};
  lineBuffer_5288 = _RAND_5295[7:0];
  _RAND_5296 = {1{`RANDOM}};
  lineBuffer_5289 = _RAND_5296[7:0];
  _RAND_5297 = {1{`RANDOM}};
  lineBuffer_5290 = _RAND_5297[7:0];
  _RAND_5298 = {1{`RANDOM}};
  lineBuffer_5291 = _RAND_5298[7:0];
  _RAND_5299 = {1{`RANDOM}};
  lineBuffer_5292 = _RAND_5299[7:0];
  _RAND_5300 = {1{`RANDOM}};
  lineBuffer_5293 = _RAND_5300[7:0];
  _RAND_5301 = {1{`RANDOM}};
  lineBuffer_5294 = _RAND_5301[7:0];
  _RAND_5302 = {1{`RANDOM}};
  lineBuffer_5295 = _RAND_5302[7:0];
  _RAND_5303 = {1{`RANDOM}};
  lineBuffer_5296 = _RAND_5303[7:0];
  _RAND_5304 = {1{`RANDOM}};
  lineBuffer_5297 = _RAND_5304[7:0];
  _RAND_5305 = {1{`RANDOM}};
  lineBuffer_5298 = _RAND_5305[7:0];
  _RAND_5306 = {1{`RANDOM}};
  lineBuffer_5299 = _RAND_5306[7:0];
  _RAND_5307 = {1{`RANDOM}};
  lineBuffer_5300 = _RAND_5307[7:0];
  _RAND_5308 = {1{`RANDOM}};
  lineBuffer_5301 = _RAND_5308[7:0];
  _RAND_5309 = {1{`RANDOM}};
  lineBuffer_5302 = _RAND_5309[7:0];
  _RAND_5310 = {1{`RANDOM}};
  lineBuffer_5303 = _RAND_5310[7:0];
  _RAND_5311 = {1{`RANDOM}};
  lineBuffer_5304 = _RAND_5311[7:0];
  _RAND_5312 = {1{`RANDOM}};
  lineBuffer_5305 = _RAND_5312[7:0];
  _RAND_5313 = {1{`RANDOM}};
  lineBuffer_5306 = _RAND_5313[7:0];
  _RAND_5314 = {1{`RANDOM}};
  lineBuffer_5307 = _RAND_5314[7:0];
  _RAND_5315 = {1{`RANDOM}};
  lineBuffer_5308 = _RAND_5315[7:0];
  _RAND_5316 = {1{`RANDOM}};
  lineBuffer_5309 = _RAND_5316[7:0];
  _RAND_5317 = {1{`RANDOM}};
  lineBuffer_5310 = _RAND_5317[7:0];
  _RAND_5318 = {1{`RANDOM}};
  lineBuffer_5311 = _RAND_5318[7:0];
  _RAND_5319 = {1{`RANDOM}};
  lineBuffer_5312 = _RAND_5319[7:0];
  _RAND_5320 = {1{`RANDOM}};
  lineBuffer_5313 = _RAND_5320[7:0];
  _RAND_5321 = {1{`RANDOM}};
  lineBuffer_5314 = _RAND_5321[7:0];
  _RAND_5322 = {1{`RANDOM}};
  lineBuffer_5315 = _RAND_5322[7:0];
  _RAND_5323 = {1{`RANDOM}};
  lineBuffer_5316 = _RAND_5323[7:0];
  _RAND_5324 = {1{`RANDOM}};
  lineBuffer_5317 = _RAND_5324[7:0];
  _RAND_5325 = {1{`RANDOM}};
  lineBuffer_5318 = _RAND_5325[7:0];
  _RAND_5326 = {1{`RANDOM}};
  lineBuffer_5319 = _RAND_5326[7:0];
  _RAND_5327 = {1{`RANDOM}};
  lineBuffer_5320 = _RAND_5327[7:0];
  _RAND_5328 = {1{`RANDOM}};
  lineBuffer_5321 = _RAND_5328[7:0];
  _RAND_5329 = {1{`RANDOM}};
  lineBuffer_5322 = _RAND_5329[7:0];
  _RAND_5330 = {1{`RANDOM}};
  lineBuffer_5323 = _RAND_5330[7:0];
  _RAND_5331 = {1{`RANDOM}};
  lineBuffer_5324 = _RAND_5331[7:0];
  _RAND_5332 = {1{`RANDOM}};
  lineBuffer_5325 = _RAND_5332[7:0];
  _RAND_5333 = {1{`RANDOM}};
  lineBuffer_5326 = _RAND_5333[7:0];
  _RAND_5334 = {1{`RANDOM}};
  lineBuffer_5327 = _RAND_5334[7:0];
  _RAND_5335 = {1{`RANDOM}};
  lineBuffer_5328 = _RAND_5335[7:0];
  _RAND_5336 = {1{`RANDOM}};
  lineBuffer_5329 = _RAND_5336[7:0];
  _RAND_5337 = {1{`RANDOM}};
  lineBuffer_5330 = _RAND_5337[7:0];
  _RAND_5338 = {1{`RANDOM}};
  lineBuffer_5331 = _RAND_5338[7:0];
  _RAND_5339 = {1{`RANDOM}};
  lineBuffer_5332 = _RAND_5339[7:0];
  _RAND_5340 = {1{`RANDOM}};
  lineBuffer_5333 = _RAND_5340[7:0];
  _RAND_5341 = {1{`RANDOM}};
  lineBuffer_5334 = _RAND_5341[7:0];
  _RAND_5342 = {1{`RANDOM}};
  lineBuffer_5335 = _RAND_5342[7:0];
  _RAND_5343 = {1{`RANDOM}};
  lineBuffer_5336 = _RAND_5343[7:0];
  _RAND_5344 = {1{`RANDOM}};
  lineBuffer_5337 = _RAND_5344[7:0];
  _RAND_5345 = {1{`RANDOM}};
  lineBuffer_5338 = _RAND_5345[7:0];
  _RAND_5346 = {1{`RANDOM}};
  lineBuffer_5339 = _RAND_5346[7:0];
  _RAND_5347 = {1{`RANDOM}};
  lineBuffer_5340 = _RAND_5347[7:0];
  _RAND_5348 = {1{`RANDOM}};
  lineBuffer_5341 = _RAND_5348[7:0];
  _RAND_5349 = {1{`RANDOM}};
  lineBuffer_5342 = _RAND_5349[7:0];
  _RAND_5350 = {1{`RANDOM}};
  lineBuffer_5343 = _RAND_5350[7:0];
  _RAND_5351 = {1{`RANDOM}};
  lineBuffer_5344 = _RAND_5351[7:0];
  _RAND_5352 = {1{`RANDOM}};
  lineBuffer_5345 = _RAND_5352[7:0];
  _RAND_5353 = {1{`RANDOM}};
  lineBuffer_5346 = _RAND_5353[7:0];
  _RAND_5354 = {1{`RANDOM}};
  lineBuffer_5347 = _RAND_5354[7:0];
  _RAND_5355 = {1{`RANDOM}};
  lineBuffer_5348 = _RAND_5355[7:0];
  _RAND_5356 = {1{`RANDOM}};
  lineBuffer_5349 = _RAND_5356[7:0];
  _RAND_5357 = {1{`RANDOM}};
  lineBuffer_5350 = _RAND_5357[7:0];
  _RAND_5358 = {1{`RANDOM}};
  lineBuffer_5351 = _RAND_5358[7:0];
  _RAND_5359 = {1{`RANDOM}};
  lineBuffer_5352 = _RAND_5359[7:0];
  _RAND_5360 = {1{`RANDOM}};
  lineBuffer_5353 = _RAND_5360[7:0];
  _RAND_5361 = {1{`RANDOM}};
  lineBuffer_5354 = _RAND_5361[7:0];
  _RAND_5362 = {1{`RANDOM}};
  lineBuffer_5355 = _RAND_5362[7:0];
  _RAND_5363 = {1{`RANDOM}};
  lineBuffer_5356 = _RAND_5363[7:0];
  _RAND_5364 = {1{`RANDOM}};
  lineBuffer_5357 = _RAND_5364[7:0];
  _RAND_5365 = {1{`RANDOM}};
  lineBuffer_5358 = _RAND_5365[7:0];
  _RAND_5366 = {1{`RANDOM}};
  lineBuffer_5359 = _RAND_5366[7:0];
  _RAND_5367 = {1{`RANDOM}};
  lineBuffer_5360 = _RAND_5367[7:0];
  _RAND_5368 = {1{`RANDOM}};
  lineBuffer_5361 = _RAND_5368[7:0];
  _RAND_5369 = {1{`RANDOM}};
  lineBuffer_5362 = _RAND_5369[7:0];
  _RAND_5370 = {1{`RANDOM}};
  lineBuffer_5363 = _RAND_5370[7:0];
  _RAND_5371 = {1{`RANDOM}};
  lineBuffer_5364 = _RAND_5371[7:0];
  _RAND_5372 = {1{`RANDOM}};
  lineBuffer_5365 = _RAND_5372[7:0];
  _RAND_5373 = {1{`RANDOM}};
  lineBuffer_5366 = _RAND_5373[7:0];
  _RAND_5374 = {1{`RANDOM}};
  lineBuffer_5367 = _RAND_5374[7:0];
  _RAND_5375 = {1{`RANDOM}};
  lineBuffer_5368 = _RAND_5375[7:0];
  _RAND_5376 = {1{`RANDOM}};
  lineBuffer_5369 = _RAND_5376[7:0];
  _RAND_5377 = {1{`RANDOM}};
  lineBuffer_5370 = _RAND_5377[7:0];
  _RAND_5378 = {1{`RANDOM}};
  lineBuffer_5371 = _RAND_5378[7:0];
  _RAND_5379 = {1{`RANDOM}};
  lineBuffer_5372 = _RAND_5379[7:0];
  _RAND_5380 = {1{`RANDOM}};
  lineBuffer_5373 = _RAND_5380[7:0];
  _RAND_5381 = {1{`RANDOM}};
  lineBuffer_5374 = _RAND_5381[7:0];
  _RAND_5382 = {1{`RANDOM}};
  lineBuffer_5375 = _RAND_5382[7:0];
  _RAND_5383 = {1{`RANDOM}};
  lineBuffer_5376 = _RAND_5383[7:0];
  _RAND_5384 = {1{`RANDOM}};
  lineBuffer_5377 = _RAND_5384[7:0];
  _RAND_5385 = {1{`RANDOM}};
  lineBuffer_5378 = _RAND_5385[7:0];
  _RAND_5386 = {1{`RANDOM}};
  lineBuffer_5379 = _RAND_5386[7:0];
  _RAND_5387 = {1{`RANDOM}};
  lineBuffer_5380 = _RAND_5387[7:0];
  _RAND_5388 = {1{`RANDOM}};
  lineBuffer_5381 = _RAND_5388[7:0];
  _RAND_5389 = {1{`RANDOM}};
  lineBuffer_5382 = _RAND_5389[7:0];
  _RAND_5390 = {1{`RANDOM}};
  lineBuffer_5383 = _RAND_5390[7:0];
  _RAND_5391 = {1{`RANDOM}};
  lineBuffer_5384 = _RAND_5391[7:0];
  _RAND_5392 = {1{`RANDOM}};
  lineBuffer_5385 = _RAND_5392[7:0];
  _RAND_5393 = {1{`RANDOM}};
  lineBuffer_5386 = _RAND_5393[7:0];
  _RAND_5394 = {1{`RANDOM}};
  lineBuffer_5387 = _RAND_5394[7:0];
  _RAND_5395 = {1{`RANDOM}};
  lineBuffer_5388 = _RAND_5395[7:0];
  _RAND_5396 = {1{`RANDOM}};
  lineBuffer_5389 = _RAND_5396[7:0];
  _RAND_5397 = {1{`RANDOM}};
  lineBuffer_5390 = _RAND_5397[7:0];
  _RAND_5398 = {1{`RANDOM}};
  lineBuffer_5391 = _RAND_5398[7:0];
  _RAND_5399 = {1{`RANDOM}};
  lineBuffer_5392 = _RAND_5399[7:0];
  _RAND_5400 = {1{`RANDOM}};
  lineBuffer_5393 = _RAND_5400[7:0];
  _RAND_5401 = {1{`RANDOM}};
  lineBuffer_5394 = _RAND_5401[7:0];
  _RAND_5402 = {1{`RANDOM}};
  lineBuffer_5395 = _RAND_5402[7:0];
  _RAND_5403 = {1{`RANDOM}};
  lineBuffer_5396 = _RAND_5403[7:0];
  _RAND_5404 = {1{`RANDOM}};
  lineBuffer_5397 = _RAND_5404[7:0];
  _RAND_5405 = {1{`RANDOM}};
  lineBuffer_5398 = _RAND_5405[7:0];
  _RAND_5406 = {1{`RANDOM}};
  lineBuffer_5399 = _RAND_5406[7:0];
  _RAND_5407 = {1{`RANDOM}};
  lineBuffer_5400 = _RAND_5407[7:0];
  _RAND_5408 = {1{`RANDOM}};
  lineBuffer_5401 = _RAND_5408[7:0];
  _RAND_5409 = {1{`RANDOM}};
  lineBuffer_5402 = _RAND_5409[7:0];
  _RAND_5410 = {1{`RANDOM}};
  lineBuffer_5403 = _RAND_5410[7:0];
  _RAND_5411 = {1{`RANDOM}};
  lineBuffer_5404 = _RAND_5411[7:0];
  _RAND_5412 = {1{`RANDOM}};
  lineBuffer_5405 = _RAND_5412[7:0];
  _RAND_5413 = {1{`RANDOM}};
  lineBuffer_5406 = _RAND_5413[7:0];
  _RAND_5414 = {1{`RANDOM}};
  lineBuffer_5407 = _RAND_5414[7:0];
  _RAND_5415 = {1{`RANDOM}};
  lineBuffer_5408 = _RAND_5415[7:0];
  _RAND_5416 = {1{`RANDOM}};
  lineBuffer_5409 = _RAND_5416[7:0];
  _RAND_5417 = {1{`RANDOM}};
  lineBuffer_5410 = _RAND_5417[7:0];
  _RAND_5418 = {1{`RANDOM}};
  lineBuffer_5411 = _RAND_5418[7:0];
  _RAND_5419 = {1{`RANDOM}};
  lineBuffer_5412 = _RAND_5419[7:0];
  _RAND_5420 = {1{`RANDOM}};
  lineBuffer_5413 = _RAND_5420[7:0];
  _RAND_5421 = {1{`RANDOM}};
  lineBuffer_5414 = _RAND_5421[7:0];
  _RAND_5422 = {1{`RANDOM}};
  lineBuffer_5415 = _RAND_5422[7:0];
  _RAND_5423 = {1{`RANDOM}};
  lineBuffer_5416 = _RAND_5423[7:0];
  _RAND_5424 = {1{`RANDOM}};
  lineBuffer_5417 = _RAND_5424[7:0];
  _RAND_5425 = {1{`RANDOM}};
  lineBuffer_5418 = _RAND_5425[7:0];
  _RAND_5426 = {1{`RANDOM}};
  lineBuffer_5419 = _RAND_5426[7:0];
  _RAND_5427 = {1{`RANDOM}};
  lineBuffer_5420 = _RAND_5427[7:0];
  _RAND_5428 = {1{`RANDOM}};
  lineBuffer_5421 = _RAND_5428[7:0];
  _RAND_5429 = {1{`RANDOM}};
  lineBuffer_5422 = _RAND_5429[7:0];
  _RAND_5430 = {1{`RANDOM}};
  lineBuffer_5423 = _RAND_5430[7:0];
  _RAND_5431 = {1{`RANDOM}};
  lineBuffer_5424 = _RAND_5431[7:0];
  _RAND_5432 = {1{`RANDOM}};
  lineBuffer_5425 = _RAND_5432[7:0];
  _RAND_5433 = {1{`RANDOM}};
  lineBuffer_5426 = _RAND_5433[7:0];
  _RAND_5434 = {1{`RANDOM}};
  lineBuffer_5427 = _RAND_5434[7:0];
  _RAND_5435 = {1{`RANDOM}};
  lineBuffer_5428 = _RAND_5435[7:0];
  _RAND_5436 = {1{`RANDOM}};
  lineBuffer_5429 = _RAND_5436[7:0];
  _RAND_5437 = {1{`RANDOM}};
  lineBuffer_5430 = _RAND_5437[7:0];
  _RAND_5438 = {1{`RANDOM}};
  lineBuffer_5431 = _RAND_5438[7:0];
  _RAND_5439 = {1{`RANDOM}};
  lineBuffer_5432 = _RAND_5439[7:0];
  _RAND_5440 = {1{`RANDOM}};
  lineBuffer_5433 = _RAND_5440[7:0];
  _RAND_5441 = {1{`RANDOM}};
  lineBuffer_5434 = _RAND_5441[7:0];
  _RAND_5442 = {1{`RANDOM}};
  lineBuffer_5435 = _RAND_5442[7:0];
  _RAND_5443 = {1{`RANDOM}};
  lineBuffer_5436 = _RAND_5443[7:0];
  _RAND_5444 = {1{`RANDOM}};
  lineBuffer_5437 = _RAND_5444[7:0];
  _RAND_5445 = {1{`RANDOM}};
  lineBuffer_5438 = _RAND_5445[7:0];
  _RAND_5446 = {1{`RANDOM}};
  lineBuffer_5439 = _RAND_5446[7:0];
  _RAND_5447 = {1{`RANDOM}};
  lineBuffer_5440 = _RAND_5447[7:0];
  _RAND_5448 = {1{`RANDOM}};
  lineBuffer_5441 = _RAND_5448[7:0];
  _RAND_5449 = {1{`RANDOM}};
  lineBuffer_5442 = _RAND_5449[7:0];
  _RAND_5450 = {1{`RANDOM}};
  lineBuffer_5443 = _RAND_5450[7:0];
  _RAND_5451 = {1{`RANDOM}};
  lineBuffer_5444 = _RAND_5451[7:0];
  _RAND_5452 = {1{`RANDOM}};
  lineBuffer_5445 = _RAND_5452[7:0];
  _RAND_5453 = {1{`RANDOM}};
  lineBuffer_5446 = _RAND_5453[7:0];
  _RAND_5454 = {1{`RANDOM}};
  lineBuffer_5447 = _RAND_5454[7:0];
  _RAND_5455 = {1{`RANDOM}};
  lineBuffer_5448 = _RAND_5455[7:0];
  _RAND_5456 = {1{`RANDOM}};
  lineBuffer_5449 = _RAND_5456[7:0];
  _RAND_5457 = {1{`RANDOM}};
  lineBuffer_5450 = _RAND_5457[7:0];
  _RAND_5458 = {1{`RANDOM}};
  lineBuffer_5451 = _RAND_5458[7:0];
  _RAND_5459 = {1{`RANDOM}};
  lineBuffer_5452 = _RAND_5459[7:0];
  _RAND_5460 = {1{`RANDOM}};
  lineBuffer_5453 = _RAND_5460[7:0];
  _RAND_5461 = {1{`RANDOM}};
  lineBuffer_5454 = _RAND_5461[7:0];
  _RAND_5462 = {1{`RANDOM}};
  lineBuffer_5455 = _RAND_5462[7:0];
  _RAND_5463 = {1{`RANDOM}};
  lineBuffer_5456 = _RAND_5463[7:0];
  _RAND_5464 = {1{`RANDOM}};
  lineBuffer_5457 = _RAND_5464[7:0];
  _RAND_5465 = {1{`RANDOM}};
  lineBuffer_5458 = _RAND_5465[7:0];
  _RAND_5466 = {1{`RANDOM}};
  lineBuffer_5459 = _RAND_5466[7:0];
  _RAND_5467 = {1{`RANDOM}};
  lineBuffer_5460 = _RAND_5467[7:0];
  _RAND_5468 = {1{`RANDOM}};
  lineBuffer_5461 = _RAND_5468[7:0];
  _RAND_5469 = {1{`RANDOM}};
  lineBuffer_5462 = _RAND_5469[7:0];
  _RAND_5470 = {1{`RANDOM}};
  lineBuffer_5463 = _RAND_5470[7:0];
  _RAND_5471 = {1{`RANDOM}};
  lineBuffer_5464 = _RAND_5471[7:0];
  _RAND_5472 = {1{`RANDOM}};
  lineBuffer_5465 = _RAND_5472[7:0];
  _RAND_5473 = {1{`RANDOM}};
  lineBuffer_5466 = _RAND_5473[7:0];
  _RAND_5474 = {1{`RANDOM}};
  lineBuffer_5467 = _RAND_5474[7:0];
  _RAND_5475 = {1{`RANDOM}};
  lineBuffer_5468 = _RAND_5475[7:0];
  _RAND_5476 = {1{`RANDOM}};
  lineBuffer_5469 = _RAND_5476[7:0];
  _RAND_5477 = {1{`RANDOM}};
  lineBuffer_5470 = _RAND_5477[7:0];
  _RAND_5478 = {1{`RANDOM}};
  lineBuffer_5471 = _RAND_5478[7:0];
  _RAND_5479 = {1{`RANDOM}};
  lineBuffer_5472 = _RAND_5479[7:0];
  _RAND_5480 = {1{`RANDOM}};
  lineBuffer_5473 = _RAND_5480[7:0];
  _RAND_5481 = {1{`RANDOM}};
  lineBuffer_5474 = _RAND_5481[7:0];
  _RAND_5482 = {1{`RANDOM}};
  lineBuffer_5475 = _RAND_5482[7:0];
  _RAND_5483 = {1{`RANDOM}};
  lineBuffer_5476 = _RAND_5483[7:0];
  _RAND_5484 = {1{`RANDOM}};
  lineBuffer_5477 = _RAND_5484[7:0];
  _RAND_5485 = {1{`RANDOM}};
  lineBuffer_5478 = _RAND_5485[7:0];
  _RAND_5486 = {1{`RANDOM}};
  lineBuffer_5479 = _RAND_5486[7:0];
  _RAND_5487 = {1{`RANDOM}};
  lineBuffer_5480 = _RAND_5487[7:0];
  _RAND_5488 = {1{`RANDOM}};
  lineBuffer_5481 = _RAND_5488[7:0];
  _RAND_5489 = {1{`RANDOM}};
  lineBuffer_5482 = _RAND_5489[7:0];
  _RAND_5490 = {1{`RANDOM}};
  lineBuffer_5483 = _RAND_5490[7:0];
  _RAND_5491 = {1{`RANDOM}};
  lineBuffer_5484 = _RAND_5491[7:0];
  _RAND_5492 = {1{`RANDOM}};
  lineBuffer_5485 = _RAND_5492[7:0];
  _RAND_5493 = {1{`RANDOM}};
  lineBuffer_5486 = _RAND_5493[7:0];
  _RAND_5494 = {1{`RANDOM}};
  lineBuffer_5487 = _RAND_5494[7:0];
  _RAND_5495 = {1{`RANDOM}};
  lineBuffer_5488 = _RAND_5495[7:0];
  _RAND_5496 = {1{`RANDOM}};
  lineBuffer_5489 = _RAND_5496[7:0];
  _RAND_5497 = {1{`RANDOM}};
  lineBuffer_5490 = _RAND_5497[7:0];
  _RAND_5498 = {1{`RANDOM}};
  lineBuffer_5491 = _RAND_5498[7:0];
  _RAND_5499 = {1{`RANDOM}};
  lineBuffer_5492 = _RAND_5499[7:0];
  _RAND_5500 = {1{`RANDOM}};
  lineBuffer_5493 = _RAND_5500[7:0];
  _RAND_5501 = {1{`RANDOM}};
  lineBuffer_5494 = _RAND_5501[7:0];
  _RAND_5502 = {1{`RANDOM}};
  lineBuffer_5495 = _RAND_5502[7:0];
  _RAND_5503 = {1{`RANDOM}};
  lineBuffer_5496 = _RAND_5503[7:0];
  _RAND_5504 = {1{`RANDOM}};
  lineBuffer_5497 = _RAND_5504[7:0];
  _RAND_5505 = {1{`RANDOM}};
  lineBuffer_5498 = _RAND_5505[7:0];
  _RAND_5506 = {1{`RANDOM}};
  lineBuffer_5499 = _RAND_5506[7:0];
  _RAND_5507 = {1{`RANDOM}};
  lineBuffer_5500 = _RAND_5507[7:0];
  _RAND_5508 = {1{`RANDOM}};
  lineBuffer_5501 = _RAND_5508[7:0];
  _RAND_5509 = {1{`RANDOM}};
  lineBuffer_5502 = _RAND_5509[7:0];
  _RAND_5510 = {1{`RANDOM}};
  lineBuffer_5503 = _RAND_5510[7:0];
  _RAND_5511 = {1{`RANDOM}};
  lineBuffer_5504 = _RAND_5511[7:0];
  _RAND_5512 = {1{`RANDOM}};
  lineBuffer_5505 = _RAND_5512[7:0];
  _RAND_5513 = {1{`RANDOM}};
  lineBuffer_5506 = _RAND_5513[7:0];
  _RAND_5514 = {1{`RANDOM}};
  lineBuffer_5507 = _RAND_5514[7:0];
  _RAND_5515 = {1{`RANDOM}};
  lineBuffer_5508 = _RAND_5515[7:0];
  _RAND_5516 = {1{`RANDOM}};
  lineBuffer_5509 = _RAND_5516[7:0];
  _RAND_5517 = {1{`RANDOM}};
  lineBuffer_5510 = _RAND_5517[7:0];
  _RAND_5518 = {1{`RANDOM}};
  lineBuffer_5511 = _RAND_5518[7:0];
  _RAND_5519 = {1{`RANDOM}};
  lineBuffer_5512 = _RAND_5519[7:0];
  _RAND_5520 = {1{`RANDOM}};
  lineBuffer_5513 = _RAND_5520[7:0];
  _RAND_5521 = {1{`RANDOM}};
  lineBuffer_5514 = _RAND_5521[7:0];
  _RAND_5522 = {1{`RANDOM}};
  lineBuffer_5515 = _RAND_5522[7:0];
  _RAND_5523 = {1{`RANDOM}};
  lineBuffer_5516 = _RAND_5523[7:0];
  _RAND_5524 = {1{`RANDOM}};
  lineBuffer_5517 = _RAND_5524[7:0];
  _RAND_5525 = {1{`RANDOM}};
  lineBuffer_5518 = _RAND_5525[7:0];
  _RAND_5526 = {1{`RANDOM}};
  lineBuffer_5519 = _RAND_5526[7:0];
  _RAND_5527 = {1{`RANDOM}};
  lineBuffer_5520 = _RAND_5527[7:0];
  _RAND_5528 = {1{`RANDOM}};
  lineBuffer_5521 = _RAND_5528[7:0];
  _RAND_5529 = {1{`RANDOM}};
  lineBuffer_5522 = _RAND_5529[7:0];
  _RAND_5530 = {1{`RANDOM}};
  lineBuffer_5523 = _RAND_5530[7:0];
  _RAND_5531 = {1{`RANDOM}};
  lineBuffer_5524 = _RAND_5531[7:0];
  _RAND_5532 = {1{`RANDOM}};
  lineBuffer_5525 = _RAND_5532[7:0];
  _RAND_5533 = {1{`RANDOM}};
  lineBuffer_5526 = _RAND_5533[7:0];
  _RAND_5534 = {1{`RANDOM}};
  lineBuffer_5527 = _RAND_5534[7:0];
  _RAND_5535 = {1{`RANDOM}};
  lineBuffer_5528 = _RAND_5535[7:0];
  _RAND_5536 = {1{`RANDOM}};
  lineBuffer_5529 = _RAND_5536[7:0];
  _RAND_5537 = {1{`RANDOM}};
  lineBuffer_5530 = _RAND_5537[7:0];
  _RAND_5538 = {1{`RANDOM}};
  lineBuffer_5531 = _RAND_5538[7:0];
  _RAND_5539 = {1{`RANDOM}};
  lineBuffer_5532 = _RAND_5539[7:0];
  _RAND_5540 = {1{`RANDOM}};
  lineBuffer_5533 = _RAND_5540[7:0];
  _RAND_5541 = {1{`RANDOM}};
  lineBuffer_5534 = _RAND_5541[7:0];
  _RAND_5542 = {1{`RANDOM}};
  lineBuffer_5535 = _RAND_5542[7:0];
  _RAND_5543 = {1{`RANDOM}};
  lineBuffer_5536 = _RAND_5543[7:0];
  _RAND_5544 = {1{`RANDOM}};
  lineBuffer_5537 = _RAND_5544[7:0];
  _RAND_5545 = {1{`RANDOM}};
  lineBuffer_5538 = _RAND_5545[7:0];
  _RAND_5546 = {1{`RANDOM}};
  lineBuffer_5539 = _RAND_5546[7:0];
  _RAND_5547 = {1{`RANDOM}};
  lineBuffer_5540 = _RAND_5547[7:0];
  _RAND_5548 = {1{`RANDOM}};
  lineBuffer_5541 = _RAND_5548[7:0];
  _RAND_5549 = {1{`RANDOM}};
  lineBuffer_5542 = _RAND_5549[7:0];
  _RAND_5550 = {1{`RANDOM}};
  lineBuffer_5543 = _RAND_5550[7:0];
  _RAND_5551 = {1{`RANDOM}};
  lineBuffer_5544 = _RAND_5551[7:0];
  _RAND_5552 = {1{`RANDOM}};
  lineBuffer_5545 = _RAND_5552[7:0];
  _RAND_5553 = {1{`RANDOM}};
  lineBuffer_5546 = _RAND_5553[7:0];
  _RAND_5554 = {1{`RANDOM}};
  lineBuffer_5547 = _RAND_5554[7:0];
  _RAND_5555 = {1{`RANDOM}};
  lineBuffer_5548 = _RAND_5555[7:0];
  _RAND_5556 = {1{`RANDOM}};
  lineBuffer_5549 = _RAND_5556[7:0];
  _RAND_5557 = {1{`RANDOM}};
  lineBuffer_5550 = _RAND_5557[7:0];
  _RAND_5558 = {1{`RANDOM}};
  lineBuffer_5551 = _RAND_5558[7:0];
  _RAND_5559 = {1{`RANDOM}};
  lineBuffer_5552 = _RAND_5559[7:0];
  _RAND_5560 = {1{`RANDOM}};
  lineBuffer_5553 = _RAND_5560[7:0];
  _RAND_5561 = {1{`RANDOM}};
  lineBuffer_5554 = _RAND_5561[7:0];
  _RAND_5562 = {1{`RANDOM}};
  lineBuffer_5555 = _RAND_5562[7:0];
  _RAND_5563 = {1{`RANDOM}};
  lineBuffer_5556 = _RAND_5563[7:0];
  _RAND_5564 = {1{`RANDOM}};
  lineBuffer_5557 = _RAND_5564[7:0];
  _RAND_5565 = {1{`RANDOM}};
  lineBuffer_5558 = _RAND_5565[7:0];
  _RAND_5566 = {1{`RANDOM}};
  lineBuffer_5559 = _RAND_5566[7:0];
  _RAND_5567 = {1{`RANDOM}};
  lineBuffer_5560 = _RAND_5567[7:0];
  _RAND_5568 = {1{`RANDOM}};
  lineBuffer_5561 = _RAND_5568[7:0];
  _RAND_5569 = {1{`RANDOM}};
  lineBuffer_5562 = _RAND_5569[7:0];
  _RAND_5570 = {1{`RANDOM}};
  lineBuffer_5563 = _RAND_5570[7:0];
  _RAND_5571 = {1{`RANDOM}};
  lineBuffer_5564 = _RAND_5571[7:0];
  _RAND_5572 = {1{`RANDOM}};
  lineBuffer_5565 = _RAND_5572[7:0];
  _RAND_5573 = {1{`RANDOM}};
  lineBuffer_5566 = _RAND_5573[7:0];
  _RAND_5574 = {1{`RANDOM}};
  lineBuffer_5567 = _RAND_5574[7:0];
  _RAND_5575 = {1{`RANDOM}};
  lineBuffer_5568 = _RAND_5575[7:0];
  _RAND_5576 = {1{`RANDOM}};
  lineBuffer_5569 = _RAND_5576[7:0];
  _RAND_5577 = {1{`RANDOM}};
  lineBuffer_5570 = _RAND_5577[7:0];
  _RAND_5578 = {1{`RANDOM}};
  lineBuffer_5571 = _RAND_5578[7:0];
  _RAND_5579 = {1{`RANDOM}};
  lineBuffer_5572 = _RAND_5579[7:0];
  _RAND_5580 = {1{`RANDOM}};
  lineBuffer_5573 = _RAND_5580[7:0];
  _RAND_5581 = {1{`RANDOM}};
  lineBuffer_5574 = _RAND_5581[7:0];
  _RAND_5582 = {1{`RANDOM}};
  lineBuffer_5575 = _RAND_5582[7:0];
  _RAND_5583 = {1{`RANDOM}};
  lineBuffer_5576 = _RAND_5583[7:0];
  _RAND_5584 = {1{`RANDOM}};
  lineBuffer_5577 = _RAND_5584[7:0];
  _RAND_5585 = {1{`RANDOM}};
  lineBuffer_5578 = _RAND_5585[7:0];
  _RAND_5586 = {1{`RANDOM}};
  lineBuffer_5579 = _RAND_5586[7:0];
  _RAND_5587 = {1{`RANDOM}};
  lineBuffer_5580 = _RAND_5587[7:0];
  _RAND_5588 = {1{`RANDOM}};
  lineBuffer_5581 = _RAND_5588[7:0];
  _RAND_5589 = {1{`RANDOM}};
  lineBuffer_5582 = _RAND_5589[7:0];
  _RAND_5590 = {1{`RANDOM}};
  lineBuffer_5583 = _RAND_5590[7:0];
  _RAND_5591 = {1{`RANDOM}};
  lineBuffer_5584 = _RAND_5591[7:0];
  _RAND_5592 = {1{`RANDOM}};
  lineBuffer_5585 = _RAND_5592[7:0];
  _RAND_5593 = {1{`RANDOM}};
  lineBuffer_5586 = _RAND_5593[7:0];
  _RAND_5594 = {1{`RANDOM}};
  lineBuffer_5587 = _RAND_5594[7:0];
  _RAND_5595 = {1{`RANDOM}};
  lineBuffer_5588 = _RAND_5595[7:0];
  _RAND_5596 = {1{`RANDOM}};
  lineBuffer_5589 = _RAND_5596[7:0];
  _RAND_5597 = {1{`RANDOM}};
  lineBuffer_5590 = _RAND_5597[7:0];
  _RAND_5598 = {1{`RANDOM}};
  lineBuffer_5591 = _RAND_5598[7:0];
  _RAND_5599 = {1{`RANDOM}};
  lineBuffer_5592 = _RAND_5599[7:0];
  _RAND_5600 = {1{`RANDOM}};
  lineBuffer_5593 = _RAND_5600[7:0];
  _RAND_5601 = {1{`RANDOM}};
  lineBuffer_5594 = _RAND_5601[7:0];
  _RAND_5602 = {1{`RANDOM}};
  lineBuffer_5595 = _RAND_5602[7:0];
  _RAND_5603 = {1{`RANDOM}};
  lineBuffer_5596 = _RAND_5603[7:0];
  _RAND_5604 = {1{`RANDOM}};
  lineBuffer_5597 = _RAND_5604[7:0];
  _RAND_5605 = {1{`RANDOM}};
  lineBuffer_5598 = _RAND_5605[7:0];
  _RAND_5606 = {1{`RANDOM}};
  lineBuffer_5599 = _RAND_5606[7:0];
  _RAND_5607 = {1{`RANDOM}};
  lineBuffer_5600 = _RAND_5607[7:0];
  _RAND_5608 = {1{`RANDOM}};
  lineBuffer_5601 = _RAND_5608[7:0];
  _RAND_5609 = {1{`RANDOM}};
  lineBuffer_5602 = _RAND_5609[7:0];
  _RAND_5610 = {1{`RANDOM}};
  lineBuffer_5603 = _RAND_5610[7:0];
  _RAND_5611 = {1{`RANDOM}};
  lineBuffer_5604 = _RAND_5611[7:0];
  _RAND_5612 = {1{`RANDOM}};
  lineBuffer_5605 = _RAND_5612[7:0];
  _RAND_5613 = {1{`RANDOM}};
  lineBuffer_5606 = _RAND_5613[7:0];
  _RAND_5614 = {1{`RANDOM}};
  lineBuffer_5607 = _RAND_5614[7:0];
  _RAND_5615 = {1{`RANDOM}};
  lineBuffer_5608 = _RAND_5615[7:0];
  _RAND_5616 = {1{`RANDOM}};
  lineBuffer_5609 = _RAND_5616[7:0];
  _RAND_5617 = {1{`RANDOM}};
  lineBuffer_5610 = _RAND_5617[7:0];
  _RAND_5618 = {1{`RANDOM}};
  lineBuffer_5611 = _RAND_5618[7:0];
  _RAND_5619 = {1{`RANDOM}};
  lineBuffer_5612 = _RAND_5619[7:0];
  _RAND_5620 = {1{`RANDOM}};
  lineBuffer_5613 = _RAND_5620[7:0];
  _RAND_5621 = {1{`RANDOM}};
  lineBuffer_5614 = _RAND_5621[7:0];
  _RAND_5622 = {1{`RANDOM}};
  lineBuffer_5615 = _RAND_5622[7:0];
  _RAND_5623 = {1{`RANDOM}};
  lineBuffer_5616 = _RAND_5623[7:0];
  _RAND_5624 = {1{`RANDOM}};
  lineBuffer_5617 = _RAND_5624[7:0];
  _RAND_5625 = {1{`RANDOM}};
  lineBuffer_5618 = _RAND_5625[7:0];
  _RAND_5626 = {1{`RANDOM}};
  lineBuffer_5619 = _RAND_5626[7:0];
  _RAND_5627 = {1{`RANDOM}};
  lineBuffer_5620 = _RAND_5627[7:0];
  _RAND_5628 = {1{`RANDOM}};
  lineBuffer_5621 = _RAND_5628[7:0];
  _RAND_5629 = {1{`RANDOM}};
  lineBuffer_5622 = _RAND_5629[7:0];
  _RAND_5630 = {1{`RANDOM}};
  lineBuffer_5623 = _RAND_5630[7:0];
  _RAND_5631 = {1{`RANDOM}};
  lineBuffer_5624 = _RAND_5631[7:0];
  _RAND_5632 = {1{`RANDOM}};
  lineBuffer_5625 = _RAND_5632[7:0];
  _RAND_5633 = {1{`RANDOM}};
  lineBuffer_5626 = _RAND_5633[7:0];
  _RAND_5634 = {1{`RANDOM}};
  lineBuffer_5627 = _RAND_5634[7:0];
  _RAND_5635 = {1{`RANDOM}};
  lineBuffer_5628 = _RAND_5635[7:0];
  _RAND_5636 = {1{`RANDOM}};
  lineBuffer_5629 = _RAND_5636[7:0];
  _RAND_5637 = {1{`RANDOM}};
  lineBuffer_5630 = _RAND_5637[7:0];
  _RAND_5638 = {1{`RANDOM}};
  lineBuffer_5631 = _RAND_5638[7:0];
  _RAND_5639 = {1{`RANDOM}};
  lineBuffer_5632 = _RAND_5639[7:0];
  _RAND_5640 = {1{`RANDOM}};
  lineBuffer_5633 = _RAND_5640[7:0];
  _RAND_5641 = {1{`RANDOM}};
  lineBuffer_5634 = _RAND_5641[7:0];
  _RAND_5642 = {1{`RANDOM}};
  lineBuffer_5635 = _RAND_5642[7:0];
  _RAND_5643 = {1{`RANDOM}};
  lineBuffer_5636 = _RAND_5643[7:0];
  _RAND_5644 = {1{`RANDOM}};
  lineBuffer_5637 = _RAND_5644[7:0];
  _RAND_5645 = {1{`RANDOM}};
  lineBuffer_5638 = _RAND_5645[7:0];
  _RAND_5646 = {1{`RANDOM}};
  lineBuffer_5639 = _RAND_5646[7:0];
  _RAND_5647 = {1{`RANDOM}};
  lineBuffer_5640 = _RAND_5647[7:0];
  _RAND_5648 = {1{`RANDOM}};
  lineBuffer_5641 = _RAND_5648[7:0];
  _RAND_5649 = {1{`RANDOM}};
  lineBuffer_5642 = _RAND_5649[7:0];
  _RAND_5650 = {1{`RANDOM}};
  lineBuffer_5643 = _RAND_5650[7:0];
  _RAND_5651 = {1{`RANDOM}};
  lineBuffer_5644 = _RAND_5651[7:0];
  _RAND_5652 = {1{`RANDOM}};
  lineBuffer_5645 = _RAND_5652[7:0];
  _RAND_5653 = {1{`RANDOM}};
  lineBuffer_5646 = _RAND_5653[7:0];
  _RAND_5654 = {1{`RANDOM}};
  lineBuffer_5647 = _RAND_5654[7:0];
  _RAND_5655 = {1{`RANDOM}};
  lineBuffer_5648 = _RAND_5655[7:0];
  _RAND_5656 = {1{`RANDOM}};
  lineBuffer_5649 = _RAND_5656[7:0];
  _RAND_5657 = {1{`RANDOM}};
  lineBuffer_5650 = _RAND_5657[7:0];
  _RAND_5658 = {1{`RANDOM}};
  lineBuffer_5651 = _RAND_5658[7:0];
  _RAND_5659 = {1{`RANDOM}};
  lineBuffer_5652 = _RAND_5659[7:0];
  _RAND_5660 = {1{`RANDOM}};
  lineBuffer_5653 = _RAND_5660[7:0];
  _RAND_5661 = {1{`RANDOM}};
  lineBuffer_5654 = _RAND_5661[7:0];
  _RAND_5662 = {1{`RANDOM}};
  lineBuffer_5655 = _RAND_5662[7:0];
  _RAND_5663 = {1{`RANDOM}};
  lineBuffer_5656 = _RAND_5663[7:0];
  _RAND_5664 = {1{`RANDOM}};
  lineBuffer_5657 = _RAND_5664[7:0];
  _RAND_5665 = {1{`RANDOM}};
  lineBuffer_5658 = _RAND_5665[7:0];
  _RAND_5666 = {1{`RANDOM}};
  lineBuffer_5659 = _RAND_5666[7:0];
  _RAND_5667 = {1{`RANDOM}};
  lineBuffer_5660 = _RAND_5667[7:0];
  _RAND_5668 = {1{`RANDOM}};
  lineBuffer_5661 = _RAND_5668[7:0];
  _RAND_5669 = {1{`RANDOM}};
  lineBuffer_5662 = _RAND_5669[7:0];
  _RAND_5670 = {1{`RANDOM}};
  lineBuffer_5663 = _RAND_5670[7:0];
  _RAND_5671 = {1{`RANDOM}};
  lineBuffer_5664 = _RAND_5671[7:0];
  _RAND_5672 = {1{`RANDOM}};
  lineBuffer_5665 = _RAND_5672[7:0];
  _RAND_5673 = {1{`RANDOM}};
  lineBuffer_5666 = _RAND_5673[7:0];
  _RAND_5674 = {1{`RANDOM}};
  lineBuffer_5667 = _RAND_5674[7:0];
  _RAND_5675 = {1{`RANDOM}};
  lineBuffer_5668 = _RAND_5675[7:0];
  _RAND_5676 = {1{`RANDOM}};
  lineBuffer_5669 = _RAND_5676[7:0];
  _RAND_5677 = {1{`RANDOM}};
  lineBuffer_5670 = _RAND_5677[7:0];
  _RAND_5678 = {1{`RANDOM}};
  lineBuffer_5671 = _RAND_5678[7:0];
  _RAND_5679 = {1{`RANDOM}};
  lineBuffer_5672 = _RAND_5679[7:0];
  _RAND_5680 = {1{`RANDOM}};
  lineBuffer_5673 = _RAND_5680[7:0];
  _RAND_5681 = {1{`RANDOM}};
  lineBuffer_5674 = _RAND_5681[7:0];
  _RAND_5682 = {1{`RANDOM}};
  lineBuffer_5675 = _RAND_5682[7:0];
  _RAND_5683 = {1{`RANDOM}};
  lineBuffer_5676 = _RAND_5683[7:0];
  _RAND_5684 = {1{`RANDOM}};
  lineBuffer_5677 = _RAND_5684[7:0];
  _RAND_5685 = {1{`RANDOM}};
  lineBuffer_5678 = _RAND_5685[7:0];
  _RAND_5686 = {1{`RANDOM}};
  lineBuffer_5679 = _RAND_5686[7:0];
  _RAND_5687 = {1{`RANDOM}};
  lineBuffer_5680 = _RAND_5687[7:0];
  _RAND_5688 = {1{`RANDOM}};
  lineBuffer_5681 = _RAND_5688[7:0];
  _RAND_5689 = {1{`RANDOM}};
  lineBuffer_5682 = _RAND_5689[7:0];
  _RAND_5690 = {1{`RANDOM}};
  lineBuffer_5683 = _RAND_5690[7:0];
  _RAND_5691 = {1{`RANDOM}};
  lineBuffer_5684 = _RAND_5691[7:0];
  _RAND_5692 = {1{`RANDOM}};
  lineBuffer_5685 = _RAND_5692[7:0];
  _RAND_5693 = {1{`RANDOM}};
  lineBuffer_5686 = _RAND_5693[7:0];
  _RAND_5694 = {1{`RANDOM}};
  lineBuffer_5687 = _RAND_5694[7:0];
  _RAND_5695 = {1{`RANDOM}};
  lineBuffer_5688 = _RAND_5695[7:0];
  _RAND_5696 = {1{`RANDOM}};
  lineBuffer_5689 = _RAND_5696[7:0];
  _RAND_5697 = {1{`RANDOM}};
  lineBuffer_5690 = _RAND_5697[7:0];
  _RAND_5698 = {1{`RANDOM}};
  lineBuffer_5691 = _RAND_5698[7:0];
  _RAND_5699 = {1{`RANDOM}};
  lineBuffer_5692 = _RAND_5699[7:0];
  _RAND_5700 = {1{`RANDOM}};
  lineBuffer_5693 = _RAND_5700[7:0];
  _RAND_5701 = {1{`RANDOM}};
  lineBuffer_5694 = _RAND_5701[7:0];
  _RAND_5702 = {1{`RANDOM}};
  lineBuffer_5695 = _RAND_5702[7:0];
  _RAND_5703 = {1{`RANDOM}};
  lineBuffer_5696 = _RAND_5703[7:0];
  _RAND_5704 = {1{`RANDOM}};
  lineBuffer_5697 = _RAND_5704[7:0];
  _RAND_5705 = {1{`RANDOM}};
  lineBuffer_5698 = _RAND_5705[7:0];
  _RAND_5706 = {1{`RANDOM}};
  lineBuffer_5699 = _RAND_5706[7:0];
  _RAND_5707 = {1{`RANDOM}};
  lineBuffer_5700 = _RAND_5707[7:0];
  _RAND_5708 = {1{`RANDOM}};
  lineBuffer_5701 = _RAND_5708[7:0];
  _RAND_5709 = {1{`RANDOM}};
  lineBuffer_5702 = _RAND_5709[7:0];
  _RAND_5710 = {1{`RANDOM}};
  lineBuffer_5703 = _RAND_5710[7:0];
  _RAND_5711 = {1{`RANDOM}};
  lineBuffer_5704 = _RAND_5711[7:0];
  _RAND_5712 = {1{`RANDOM}};
  lineBuffer_5705 = _RAND_5712[7:0];
  _RAND_5713 = {1{`RANDOM}};
  lineBuffer_5706 = _RAND_5713[7:0];
  _RAND_5714 = {1{`RANDOM}};
  lineBuffer_5707 = _RAND_5714[7:0];
  _RAND_5715 = {1{`RANDOM}};
  lineBuffer_5708 = _RAND_5715[7:0];
  _RAND_5716 = {1{`RANDOM}};
  lineBuffer_5709 = _RAND_5716[7:0];
  _RAND_5717 = {1{`RANDOM}};
  lineBuffer_5710 = _RAND_5717[7:0];
  _RAND_5718 = {1{`RANDOM}};
  lineBuffer_5711 = _RAND_5718[7:0];
  _RAND_5719 = {1{`RANDOM}};
  lineBuffer_5712 = _RAND_5719[7:0];
  _RAND_5720 = {1{`RANDOM}};
  lineBuffer_5713 = _RAND_5720[7:0];
  _RAND_5721 = {1{`RANDOM}};
  lineBuffer_5714 = _RAND_5721[7:0];
  _RAND_5722 = {1{`RANDOM}};
  lineBuffer_5715 = _RAND_5722[7:0];
  _RAND_5723 = {1{`RANDOM}};
  lineBuffer_5716 = _RAND_5723[7:0];
  _RAND_5724 = {1{`RANDOM}};
  lineBuffer_5717 = _RAND_5724[7:0];
  _RAND_5725 = {1{`RANDOM}};
  lineBuffer_5718 = _RAND_5725[7:0];
  _RAND_5726 = {1{`RANDOM}};
  lineBuffer_5719 = _RAND_5726[7:0];
  _RAND_5727 = {1{`RANDOM}};
  lineBuffer_5720 = _RAND_5727[7:0];
  _RAND_5728 = {1{`RANDOM}};
  lineBuffer_5721 = _RAND_5728[7:0];
  _RAND_5729 = {1{`RANDOM}};
  lineBuffer_5722 = _RAND_5729[7:0];
  _RAND_5730 = {1{`RANDOM}};
  lineBuffer_5723 = _RAND_5730[7:0];
  _RAND_5731 = {1{`RANDOM}};
  lineBuffer_5724 = _RAND_5731[7:0];
  _RAND_5732 = {1{`RANDOM}};
  lineBuffer_5725 = _RAND_5732[7:0];
  _RAND_5733 = {1{`RANDOM}};
  lineBuffer_5726 = _RAND_5733[7:0];
  _RAND_5734 = {1{`RANDOM}};
  lineBuffer_5727 = _RAND_5734[7:0];
  _RAND_5735 = {1{`RANDOM}};
  lineBuffer_5728 = _RAND_5735[7:0];
  _RAND_5736 = {1{`RANDOM}};
  lineBuffer_5729 = _RAND_5736[7:0];
  _RAND_5737 = {1{`RANDOM}};
  lineBuffer_5730 = _RAND_5737[7:0];
  _RAND_5738 = {1{`RANDOM}};
  lineBuffer_5731 = _RAND_5738[7:0];
  _RAND_5739 = {1{`RANDOM}};
  lineBuffer_5732 = _RAND_5739[7:0];
  _RAND_5740 = {1{`RANDOM}};
  lineBuffer_5733 = _RAND_5740[7:0];
  _RAND_5741 = {1{`RANDOM}};
  lineBuffer_5734 = _RAND_5741[7:0];
  _RAND_5742 = {1{`RANDOM}};
  lineBuffer_5735 = _RAND_5742[7:0];
  _RAND_5743 = {1{`RANDOM}};
  lineBuffer_5736 = _RAND_5743[7:0];
  _RAND_5744 = {1{`RANDOM}};
  lineBuffer_5737 = _RAND_5744[7:0];
  _RAND_5745 = {1{`RANDOM}};
  lineBuffer_5738 = _RAND_5745[7:0];
  _RAND_5746 = {1{`RANDOM}};
  lineBuffer_5739 = _RAND_5746[7:0];
  _RAND_5747 = {1{`RANDOM}};
  lineBuffer_5740 = _RAND_5747[7:0];
  _RAND_5748 = {1{`RANDOM}};
  lineBuffer_5741 = _RAND_5748[7:0];
  _RAND_5749 = {1{`RANDOM}};
  lineBuffer_5742 = _RAND_5749[7:0];
  _RAND_5750 = {1{`RANDOM}};
  lineBuffer_5743 = _RAND_5750[7:0];
  _RAND_5751 = {1{`RANDOM}};
  lineBuffer_5744 = _RAND_5751[7:0];
  _RAND_5752 = {1{`RANDOM}};
  lineBuffer_5745 = _RAND_5752[7:0];
  _RAND_5753 = {1{`RANDOM}};
  lineBuffer_5746 = _RAND_5753[7:0];
  _RAND_5754 = {1{`RANDOM}};
  lineBuffer_5747 = _RAND_5754[7:0];
  _RAND_5755 = {1{`RANDOM}};
  lineBuffer_5748 = _RAND_5755[7:0];
  _RAND_5756 = {1{`RANDOM}};
  lineBuffer_5749 = _RAND_5756[7:0];
  _RAND_5757 = {1{`RANDOM}};
  lineBuffer_5750 = _RAND_5757[7:0];
  _RAND_5758 = {1{`RANDOM}};
  lineBuffer_5751 = _RAND_5758[7:0];
  _RAND_5759 = {1{`RANDOM}};
  lineBuffer_5752 = _RAND_5759[7:0];
  _RAND_5760 = {1{`RANDOM}};
  lineBuffer_5753 = _RAND_5760[7:0];
  _RAND_5761 = {1{`RANDOM}};
  lineBuffer_5754 = _RAND_5761[7:0];
  _RAND_5762 = {1{`RANDOM}};
  lineBuffer_5755 = _RAND_5762[7:0];
  _RAND_5763 = {1{`RANDOM}};
  lineBuffer_5756 = _RAND_5763[7:0];
  _RAND_5764 = {1{`RANDOM}};
  lineBuffer_5757 = _RAND_5764[7:0];
  _RAND_5765 = {1{`RANDOM}};
  lineBuffer_5758 = _RAND_5765[7:0];
  _RAND_5766 = {1{`RANDOM}};
  lineBuffer_5759 = _RAND_5766[7:0];
  _RAND_5767 = {1{`RANDOM}};
  lineBuffer_5760 = _RAND_5767[7:0];
  _RAND_5768 = {1{`RANDOM}};
  lineBuffer_5761 = _RAND_5768[7:0];
  _RAND_5769 = {1{`RANDOM}};
  lineBuffer_5762 = _RAND_5769[7:0];
  _RAND_5770 = {1{`RANDOM}};
  lineBuffer_5763 = _RAND_5770[7:0];
  _RAND_5771 = {1{`RANDOM}};
  lineBuffer_5764 = _RAND_5771[7:0];
  _RAND_5772 = {1{`RANDOM}};
  lineBuffer_5765 = _RAND_5772[7:0];
  _RAND_5773 = {1{`RANDOM}};
  lineBuffer_5766 = _RAND_5773[7:0];
  _RAND_5774 = {1{`RANDOM}};
  lineBuffer_5767 = _RAND_5774[7:0];
  _RAND_5775 = {1{`RANDOM}};
  lineBuffer_5768 = _RAND_5775[7:0];
  _RAND_5776 = {1{`RANDOM}};
  lineBuffer_5769 = _RAND_5776[7:0];
  _RAND_5777 = {1{`RANDOM}};
  lineBuffer_5770 = _RAND_5777[7:0];
  _RAND_5778 = {1{`RANDOM}};
  lineBuffer_5771 = _RAND_5778[7:0];
  _RAND_5779 = {1{`RANDOM}};
  lineBuffer_5772 = _RAND_5779[7:0];
  _RAND_5780 = {1{`RANDOM}};
  lineBuffer_5773 = _RAND_5780[7:0];
  _RAND_5781 = {1{`RANDOM}};
  lineBuffer_5774 = _RAND_5781[7:0];
  _RAND_5782 = {1{`RANDOM}};
  lineBuffer_5775 = _RAND_5782[7:0];
  _RAND_5783 = {1{`RANDOM}};
  lineBuffer_5776 = _RAND_5783[7:0];
  _RAND_5784 = {1{`RANDOM}};
  lineBuffer_5777 = _RAND_5784[7:0];
  _RAND_5785 = {1{`RANDOM}};
  lineBuffer_5778 = _RAND_5785[7:0];
  _RAND_5786 = {1{`RANDOM}};
  lineBuffer_5779 = _RAND_5786[7:0];
  _RAND_5787 = {1{`RANDOM}};
  lineBuffer_5780 = _RAND_5787[7:0];
  _RAND_5788 = {1{`RANDOM}};
  lineBuffer_5781 = _RAND_5788[7:0];
  _RAND_5789 = {1{`RANDOM}};
  lineBuffer_5782 = _RAND_5789[7:0];
  _RAND_5790 = {1{`RANDOM}};
  lineBuffer_5783 = _RAND_5790[7:0];
  _RAND_5791 = {1{`RANDOM}};
  lineBuffer_5784 = _RAND_5791[7:0];
  _RAND_5792 = {1{`RANDOM}};
  lineBuffer_5785 = _RAND_5792[7:0];
  _RAND_5793 = {1{`RANDOM}};
  lineBuffer_5786 = _RAND_5793[7:0];
  _RAND_5794 = {1{`RANDOM}};
  lineBuffer_5787 = _RAND_5794[7:0];
  _RAND_5795 = {1{`RANDOM}};
  lineBuffer_5788 = _RAND_5795[7:0];
  _RAND_5796 = {1{`RANDOM}};
  lineBuffer_5789 = _RAND_5796[7:0];
  _RAND_5797 = {1{`RANDOM}};
  lineBuffer_5790 = _RAND_5797[7:0];
  _RAND_5798 = {1{`RANDOM}};
  lineBuffer_5791 = _RAND_5798[7:0];
  _RAND_5799 = {1{`RANDOM}};
  lineBuffer_5792 = _RAND_5799[7:0];
  _RAND_5800 = {1{`RANDOM}};
  lineBuffer_5793 = _RAND_5800[7:0];
  _RAND_5801 = {1{`RANDOM}};
  lineBuffer_5794 = _RAND_5801[7:0];
  _RAND_5802 = {1{`RANDOM}};
  lineBuffer_5795 = _RAND_5802[7:0];
  _RAND_5803 = {1{`RANDOM}};
  lineBuffer_5796 = _RAND_5803[7:0];
  _RAND_5804 = {1{`RANDOM}};
  lineBuffer_5797 = _RAND_5804[7:0];
  _RAND_5805 = {1{`RANDOM}};
  lineBuffer_5798 = _RAND_5805[7:0];
  _RAND_5806 = {1{`RANDOM}};
  lineBuffer_5799 = _RAND_5806[7:0];
  _RAND_5807 = {1{`RANDOM}};
  lineBuffer_5800 = _RAND_5807[7:0];
  _RAND_5808 = {1{`RANDOM}};
  lineBuffer_5801 = _RAND_5808[7:0];
  _RAND_5809 = {1{`RANDOM}};
  lineBuffer_5802 = _RAND_5809[7:0];
  _RAND_5810 = {1{`RANDOM}};
  lineBuffer_5803 = _RAND_5810[7:0];
  _RAND_5811 = {1{`RANDOM}};
  lineBuffer_5804 = _RAND_5811[7:0];
  _RAND_5812 = {1{`RANDOM}};
  lineBuffer_5805 = _RAND_5812[7:0];
  _RAND_5813 = {1{`RANDOM}};
  lineBuffer_5806 = _RAND_5813[7:0];
  _RAND_5814 = {1{`RANDOM}};
  lineBuffer_5807 = _RAND_5814[7:0];
  _RAND_5815 = {1{`RANDOM}};
  lineBuffer_5808 = _RAND_5815[7:0];
  _RAND_5816 = {1{`RANDOM}};
  lineBuffer_5809 = _RAND_5816[7:0];
  _RAND_5817 = {1{`RANDOM}};
  lineBuffer_5810 = _RAND_5817[7:0];
  _RAND_5818 = {1{`RANDOM}};
  lineBuffer_5811 = _RAND_5818[7:0];
  _RAND_5819 = {1{`RANDOM}};
  lineBuffer_5812 = _RAND_5819[7:0];
  _RAND_5820 = {1{`RANDOM}};
  lineBuffer_5813 = _RAND_5820[7:0];
  _RAND_5821 = {1{`RANDOM}};
  lineBuffer_5814 = _RAND_5821[7:0];
  _RAND_5822 = {1{`RANDOM}};
  lineBuffer_5815 = _RAND_5822[7:0];
  _RAND_5823 = {1{`RANDOM}};
  lineBuffer_5816 = _RAND_5823[7:0];
  _RAND_5824 = {1{`RANDOM}};
  lineBuffer_5817 = _RAND_5824[7:0];
  _RAND_5825 = {1{`RANDOM}};
  lineBuffer_5818 = _RAND_5825[7:0];
  _RAND_5826 = {1{`RANDOM}};
  lineBuffer_5819 = _RAND_5826[7:0];
  _RAND_5827 = {1{`RANDOM}};
  lineBuffer_5820 = _RAND_5827[7:0];
  _RAND_5828 = {1{`RANDOM}};
  lineBuffer_5821 = _RAND_5828[7:0];
  _RAND_5829 = {1{`RANDOM}};
  lineBuffer_5822 = _RAND_5829[7:0];
  _RAND_5830 = {1{`RANDOM}};
  lineBuffer_5823 = _RAND_5830[7:0];
  _RAND_5831 = {1{`RANDOM}};
  lineBuffer_5824 = _RAND_5831[7:0];
  _RAND_5832 = {1{`RANDOM}};
  lineBuffer_5825 = _RAND_5832[7:0];
  _RAND_5833 = {1{`RANDOM}};
  lineBuffer_5826 = _RAND_5833[7:0];
  _RAND_5834 = {1{`RANDOM}};
  lineBuffer_5827 = _RAND_5834[7:0];
  _RAND_5835 = {1{`RANDOM}};
  lineBuffer_5828 = _RAND_5835[7:0];
  _RAND_5836 = {1{`RANDOM}};
  lineBuffer_5829 = _RAND_5836[7:0];
  _RAND_5837 = {1{`RANDOM}};
  lineBuffer_5830 = _RAND_5837[7:0];
  _RAND_5838 = {1{`RANDOM}};
  lineBuffer_5831 = _RAND_5838[7:0];
  _RAND_5839 = {1{`RANDOM}};
  lineBuffer_5832 = _RAND_5839[7:0];
  _RAND_5840 = {1{`RANDOM}};
  lineBuffer_5833 = _RAND_5840[7:0];
  _RAND_5841 = {1{`RANDOM}};
  lineBuffer_5834 = _RAND_5841[7:0];
  _RAND_5842 = {1{`RANDOM}};
  lineBuffer_5835 = _RAND_5842[7:0];
  _RAND_5843 = {1{`RANDOM}};
  lineBuffer_5836 = _RAND_5843[7:0];
  _RAND_5844 = {1{`RANDOM}};
  lineBuffer_5837 = _RAND_5844[7:0];
  _RAND_5845 = {1{`RANDOM}};
  lineBuffer_5838 = _RAND_5845[7:0];
  _RAND_5846 = {1{`RANDOM}};
  lineBuffer_5839 = _RAND_5846[7:0];
  _RAND_5847 = {1{`RANDOM}};
  lineBuffer_5840 = _RAND_5847[7:0];
  _RAND_5848 = {1{`RANDOM}};
  lineBuffer_5841 = _RAND_5848[7:0];
  _RAND_5849 = {1{`RANDOM}};
  lineBuffer_5842 = _RAND_5849[7:0];
  _RAND_5850 = {1{`RANDOM}};
  lineBuffer_5843 = _RAND_5850[7:0];
  _RAND_5851 = {1{`RANDOM}};
  lineBuffer_5844 = _RAND_5851[7:0];
  _RAND_5852 = {1{`RANDOM}};
  lineBuffer_5845 = _RAND_5852[7:0];
  _RAND_5853 = {1{`RANDOM}};
  lineBuffer_5846 = _RAND_5853[7:0];
  _RAND_5854 = {1{`RANDOM}};
  lineBuffer_5847 = _RAND_5854[7:0];
  _RAND_5855 = {1{`RANDOM}};
  lineBuffer_5848 = _RAND_5855[7:0];
  _RAND_5856 = {1{`RANDOM}};
  lineBuffer_5849 = _RAND_5856[7:0];
  _RAND_5857 = {1{`RANDOM}};
  lineBuffer_5850 = _RAND_5857[7:0];
  _RAND_5858 = {1{`RANDOM}};
  lineBuffer_5851 = _RAND_5858[7:0];
  _RAND_5859 = {1{`RANDOM}};
  lineBuffer_5852 = _RAND_5859[7:0];
  _RAND_5860 = {1{`RANDOM}};
  lineBuffer_5853 = _RAND_5860[7:0];
  _RAND_5861 = {1{`RANDOM}};
  lineBuffer_5854 = _RAND_5861[7:0];
  _RAND_5862 = {1{`RANDOM}};
  lineBuffer_5855 = _RAND_5862[7:0];
  _RAND_5863 = {1{`RANDOM}};
  lineBuffer_5856 = _RAND_5863[7:0];
  _RAND_5864 = {1{`RANDOM}};
  lineBuffer_5857 = _RAND_5864[7:0];
  _RAND_5865 = {1{`RANDOM}};
  lineBuffer_5858 = _RAND_5865[7:0];
  _RAND_5866 = {1{`RANDOM}};
  lineBuffer_5859 = _RAND_5866[7:0];
  _RAND_5867 = {1{`RANDOM}};
  lineBuffer_5860 = _RAND_5867[7:0];
  _RAND_5868 = {1{`RANDOM}};
  lineBuffer_5861 = _RAND_5868[7:0];
  _RAND_5869 = {1{`RANDOM}};
  lineBuffer_5862 = _RAND_5869[7:0];
  _RAND_5870 = {1{`RANDOM}};
  lineBuffer_5863 = _RAND_5870[7:0];
  _RAND_5871 = {1{`RANDOM}};
  lineBuffer_5864 = _RAND_5871[7:0];
  _RAND_5872 = {1{`RANDOM}};
  lineBuffer_5865 = _RAND_5872[7:0];
  _RAND_5873 = {1{`RANDOM}};
  lineBuffer_5866 = _RAND_5873[7:0];
  _RAND_5874 = {1{`RANDOM}};
  lineBuffer_5867 = _RAND_5874[7:0];
  _RAND_5875 = {1{`RANDOM}};
  lineBuffer_5868 = _RAND_5875[7:0];
  _RAND_5876 = {1{`RANDOM}};
  lineBuffer_5869 = _RAND_5876[7:0];
  _RAND_5877 = {1{`RANDOM}};
  lineBuffer_5870 = _RAND_5877[7:0];
  _RAND_5878 = {1{`RANDOM}};
  lineBuffer_5871 = _RAND_5878[7:0];
  _RAND_5879 = {1{`RANDOM}};
  lineBuffer_5872 = _RAND_5879[7:0];
  _RAND_5880 = {1{`RANDOM}};
  lineBuffer_5873 = _RAND_5880[7:0];
  _RAND_5881 = {1{`RANDOM}};
  lineBuffer_5874 = _RAND_5881[7:0];
  _RAND_5882 = {1{`RANDOM}};
  lineBuffer_5875 = _RAND_5882[7:0];
  _RAND_5883 = {1{`RANDOM}};
  lineBuffer_5876 = _RAND_5883[7:0];
  _RAND_5884 = {1{`RANDOM}};
  lineBuffer_5877 = _RAND_5884[7:0];
  _RAND_5885 = {1{`RANDOM}};
  lineBuffer_5878 = _RAND_5885[7:0];
  _RAND_5886 = {1{`RANDOM}};
  lineBuffer_5879 = _RAND_5886[7:0];
  _RAND_5887 = {1{`RANDOM}};
  lineBuffer_5880 = _RAND_5887[7:0];
  _RAND_5888 = {1{`RANDOM}};
  lineBuffer_5881 = _RAND_5888[7:0];
  _RAND_5889 = {1{`RANDOM}};
  lineBuffer_5882 = _RAND_5889[7:0];
  _RAND_5890 = {1{`RANDOM}};
  lineBuffer_5883 = _RAND_5890[7:0];
  _RAND_5891 = {1{`RANDOM}};
  lineBuffer_5884 = _RAND_5891[7:0];
  _RAND_5892 = {1{`RANDOM}};
  lineBuffer_5885 = _RAND_5892[7:0];
  _RAND_5893 = {1{`RANDOM}};
  lineBuffer_5886 = _RAND_5893[7:0];
  _RAND_5894 = {1{`RANDOM}};
  lineBuffer_5887 = _RAND_5894[7:0];
  _RAND_5895 = {1{`RANDOM}};
  lineBuffer_5888 = _RAND_5895[7:0];
  _RAND_5896 = {1{`RANDOM}};
  lineBuffer_5889 = _RAND_5896[7:0];
  _RAND_5897 = {1{`RANDOM}};
  lineBuffer_5890 = _RAND_5897[7:0];
  _RAND_5898 = {1{`RANDOM}};
  lineBuffer_5891 = _RAND_5898[7:0];
  _RAND_5899 = {1{`RANDOM}};
  lineBuffer_5892 = _RAND_5899[7:0];
  _RAND_5900 = {1{`RANDOM}};
  lineBuffer_5893 = _RAND_5900[7:0];
  _RAND_5901 = {1{`RANDOM}};
  lineBuffer_5894 = _RAND_5901[7:0];
  _RAND_5902 = {1{`RANDOM}};
  lineBuffer_5895 = _RAND_5902[7:0];
  _RAND_5903 = {1{`RANDOM}};
  lineBuffer_5896 = _RAND_5903[7:0];
  _RAND_5904 = {1{`RANDOM}};
  lineBuffer_5897 = _RAND_5904[7:0];
  _RAND_5905 = {1{`RANDOM}};
  lineBuffer_5898 = _RAND_5905[7:0];
  _RAND_5906 = {1{`RANDOM}};
  lineBuffer_5899 = _RAND_5906[7:0];
  _RAND_5907 = {1{`RANDOM}};
  lineBuffer_5900 = _RAND_5907[7:0];
  _RAND_5908 = {1{`RANDOM}};
  lineBuffer_5901 = _RAND_5908[7:0];
  _RAND_5909 = {1{`RANDOM}};
  lineBuffer_5902 = _RAND_5909[7:0];
  _RAND_5910 = {1{`RANDOM}};
  lineBuffer_5903 = _RAND_5910[7:0];
  _RAND_5911 = {1{`RANDOM}};
  lineBuffer_5904 = _RAND_5911[7:0];
  _RAND_5912 = {1{`RANDOM}};
  lineBuffer_5905 = _RAND_5912[7:0];
  _RAND_5913 = {1{`RANDOM}};
  lineBuffer_5906 = _RAND_5913[7:0];
  _RAND_5914 = {1{`RANDOM}};
  lineBuffer_5907 = _RAND_5914[7:0];
  _RAND_5915 = {1{`RANDOM}};
  lineBuffer_5908 = _RAND_5915[7:0];
  _RAND_5916 = {1{`RANDOM}};
  lineBuffer_5909 = _RAND_5916[7:0];
  _RAND_5917 = {1{`RANDOM}};
  lineBuffer_5910 = _RAND_5917[7:0];
  _RAND_5918 = {1{`RANDOM}};
  lineBuffer_5911 = _RAND_5918[7:0];
  _RAND_5919 = {1{`RANDOM}};
  lineBuffer_5912 = _RAND_5919[7:0];
  _RAND_5920 = {1{`RANDOM}};
  lineBuffer_5913 = _RAND_5920[7:0];
  _RAND_5921 = {1{`RANDOM}};
  lineBuffer_5914 = _RAND_5921[7:0];
  _RAND_5922 = {1{`RANDOM}};
  lineBuffer_5915 = _RAND_5922[7:0];
  _RAND_5923 = {1{`RANDOM}};
  lineBuffer_5916 = _RAND_5923[7:0];
  _RAND_5924 = {1{`RANDOM}};
  lineBuffer_5917 = _RAND_5924[7:0];
  _RAND_5925 = {1{`RANDOM}};
  lineBuffer_5918 = _RAND_5925[7:0];
  _RAND_5926 = {1{`RANDOM}};
  lineBuffer_5919 = _RAND_5926[7:0];
  _RAND_5927 = {1{`RANDOM}};
  lineBuffer_5920 = _RAND_5927[7:0];
  _RAND_5928 = {1{`RANDOM}};
  lineBuffer_5921 = _RAND_5928[7:0];
  _RAND_5929 = {1{`RANDOM}};
  lineBuffer_5922 = _RAND_5929[7:0];
  _RAND_5930 = {1{`RANDOM}};
  lineBuffer_5923 = _RAND_5930[7:0];
  _RAND_5931 = {1{`RANDOM}};
  lineBuffer_5924 = _RAND_5931[7:0];
  _RAND_5932 = {1{`RANDOM}};
  lineBuffer_5925 = _RAND_5932[7:0];
  _RAND_5933 = {1{`RANDOM}};
  lineBuffer_5926 = _RAND_5933[7:0];
  _RAND_5934 = {1{`RANDOM}};
  lineBuffer_5927 = _RAND_5934[7:0];
  _RAND_5935 = {1{`RANDOM}};
  lineBuffer_5928 = _RAND_5935[7:0];
  _RAND_5936 = {1{`RANDOM}};
  lineBuffer_5929 = _RAND_5936[7:0];
  _RAND_5937 = {1{`RANDOM}};
  lineBuffer_5930 = _RAND_5937[7:0];
  _RAND_5938 = {1{`RANDOM}};
  lineBuffer_5931 = _RAND_5938[7:0];
  _RAND_5939 = {1{`RANDOM}};
  lineBuffer_5932 = _RAND_5939[7:0];
  _RAND_5940 = {1{`RANDOM}};
  lineBuffer_5933 = _RAND_5940[7:0];
  _RAND_5941 = {1{`RANDOM}};
  lineBuffer_5934 = _RAND_5941[7:0];
  _RAND_5942 = {1{`RANDOM}};
  lineBuffer_5935 = _RAND_5942[7:0];
  _RAND_5943 = {1{`RANDOM}};
  lineBuffer_5936 = _RAND_5943[7:0];
  _RAND_5944 = {1{`RANDOM}};
  lineBuffer_5937 = _RAND_5944[7:0];
  _RAND_5945 = {1{`RANDOM}};
  lineBuffer_5938 = _RAND_5945[7:0];
  _RAND_5946 = {1{`RANDOM}};
  lineBuffer_5939 = _RAND_5946[7:0];
  _RAND_5947 = {1{`RANDOM}};
  lineBuffer_5940 = _RAND_5947[7:0];
  _RAND_5948 = {1{`RANDOM}};
  lineBuffer_5941 = _RAND_5948[7:0];
  _RAND_5949 = {1{`RANDOM}};
  lineBuffer_5942 = _RAND_5949[7:0];
  _RAND_5950 = {1{`RANDOM}};
  lineBuffer_5943 = _RAND_5950[7:0];
  _RAND_5951 = {1{`RANDOM}};
  lineBuffer_5944 = _RAND_5951[7:0];
  _RAND_5952 = {1{`RANDOM}};
  lineBuffer_5945 = _RAND_5952[7:0];
  _RAND_5953 = {1{`RANDOM}};
  lineBuffer_5946 = _RAND_5953[7:0];
  _RAND_5954 = {1{`RANDOM}};
  lineBuffer_5947 = _RAND_5954[7:0];
  _RAND_5955 = {1{`RANDOM}};
  lineBuffer_5948 = _RAND_5955[7:0];
  _RAND_5956 = {1{`RANDOM}};
  lineBuffer_5949 = _RAND_5956[7:0];
  _RAND_5957 = {1{`RANDOM}};
  lineBuffer_5950 = _RAND_5957[7:0];
  _RAND_5958 = {1{`RANDOM}};
  lineBuffer_5951 = _RAND_5958[7:0];
  _RAND_5959 = {1{`RANDOM}};
  lineBuffer_5952 = _RAND_5959[7:0];
  _RAND_5960 = {1{`RANDOM}};
  lineBuffer_5953 = _RAND_5960[7:0];
  _RAND_5961 = {1{`RANDOM}};
  lineBuffer_5954 = _RAND_5961[7:0];
  _RAND_5962 = {1{`RANDOM}};
  lineBuffer_5955 = _RAND_5962[7:0];
  _RAND_5963 = {1{`RANDOM}};
  lineBuffer_5956 = _RAND_5963[7:0];
  _RAND_5964 = {1{`RANDOM}};
  lineBuffer_5957 = _RAND_5964[7:0];
  _RAND_5965 = {1{`RANDOM}};
  lineBuffer_5958 = _RAND_5965[7:0];
  _RAND_5966 = {1{`RANDOM}};
  lineBuffer_5959 = _RAND_5966[7:0];
  _RAND_5967 = {1{`RANDOM}};
  lineBuffer_5960 = _RAND_5967[7:0];
  _RAND_5968 = {1{`RANDOM}};
  lineBuffer_5961 = _RAND_5968[7:0];
  _RAND_5969 = {1{`RANDOM}};
  lineBuffer_5962 = _RAND_5969[7:0];
  _RAND_5970 = {1{`RANDOM}};
  lineBuffer_5963 = _RAND_5970[7:0];
  _RAND_5971 = {1{`RANDOM}};
  lineBuffer_5964 = _RAND_5971[7:0];
  _RAND_5972 = {1{`RANDOM}};
  lineBuffer_5965 = _RAND_5972[7:0];
  _RAND_5973 = {1{`RANDOM}};
  lineBuffer_5966 = _RAND_5973[7:0];
  _RAND_5974 = {1{`RANDOM}};
  lineBuffer_5967 = _RAND_5974[7:0];
  _RAND_5975 = {1{`RANDOM}};
  lineBuffer_5968 = _RAND_5975[7:0];
  _RAND_5976 = {1{`RANDOM}};
  lineBuffer_5969 = _RAND_5976[7:0];
  _RAND_5977 = {1{`RANDOM}};
  lineBuffer_5970 = _RAND_5977[7:0];
  _RAND_5978 = {1{`RANDOM}};
  lineBuffer_5971 = _RAND_5978[7:0];
  _RAND_5979 = {1{`RANDOM}};
  lineBuffer_5972 = _RAND_5979[7:0];
  _RAND_5980 = {1{`RANDOM}};
  lineBuffer_5973 = _RAND_5980[7:0];
  _RAND_5981 = {1{`RANDOM}};
  lineBuffer_5974 = _RAND_5981[7:0];
  _RAND_5982 = {1{`RANDOM}};
  lineBuffer_5975 = _RAND_5982[7:0];
  _RAND_5983 = {1{`RANDOM}};
  lineBuffer_5976 = _RAND_5983[7:0];
  _RAND_5984 = {1{`RANDOM}};
  lineBuffer_5977 = _RAND_5984[7:0];
  _RAND_5985 = {1{`RANDOM}};
  lineBuffer_5978 = _RAND_5985[7:0];
  _RAND_5986 = {1{`RANDOM}};
  lineBuffer_5979 = _RAND_5986[7:0];
  _RAND_5987 = {1{`RANDOM}};
  lineBuffer_5980 = _RAND_5987[7:0];
  _RAND_5988 = {1{`RANDOM}};
  lineBuffer_5981 = _RAND_5988[7:0];
  _RAND_5989 = {1{`RANDOM}};
  lineBuffer_5982 = _RAND_5989[7:0];
  _RAND_5990 = {1{`RANDOM}};
  lineBuffer_5983 = _RAND_5990[7:0];
  _RAND_5991 = {1{`RANDOM}};
  lineBuffer_5984 = _RAND_5991[7:0];
  _RAND_5992 = {1{`RANDOM}};
  lineBuffer_5985 = _RAND_5992[7:0];
  _RAND_5993 = {1{`RANDOM}};
  lineBuffer_5986 = _RAND_5993[7:0];
  _RAND_5994 = {1{`RANDOM}};
  lineBuffer_5987 = _RAND_5994[7:0];
  _RAND_5995 = {1{`RANDOM}};
  lineBuffer_5988 = _RAND_5995[7:0];
  _RAND_5996 = {1{`RANDOM}};
  lineBuffer_5989 = _RAND_5996[7:0];
  _RAND_5997 = {1{`RANDOM}};
  lineBuffer_5990 = _RAND_5997[7:0];
  _RAND_5998 = {1{`RANDOM}};
  lineBuffer_5991 = _RAND_5998[7:0];
  _RAND_5999 = {1{`RANDOM}};
  lineBuffer_5992 = _RAND_5999[7:0];
  _RAND_6000 = {1{`RANDOM}};
  lineBuffer_5993 = _RAND_6000[7:0];
  _RAND_6001 = {1{`RANDOM}};
  lineBuffer_5994 = _RAND_6001[7:0];
  _RAND_6002 = {1{`RANDOM}};
  lineBuffer_5995 = _RAND_6002[7:0];
  _RAND_6003 = {1{`RANDOM}};
  lineBuffer_5996 = _RAND_6003[7:0];
  _RAND_6004 = {1{`RANDOM}};
  lineBuffer_5997 = _RAND_6004[7:0];
  _RAND_6005 = {1{`RANDOM}};
  lineBuffer_5998 = _RAND_6005[7:0];
  _RAND_6006 = {1{`RANDOM}};
  lineBuffer_5999 = _RAND_6006[7:0];
  _RAND_6007 = {1{`RANDOM}};
  lineBuffer_6000 = _RAND_6007[7:0];
  _RAND_6008 = {1{`RANDOM}};
  lineBuffer_6001 = _RAND_6008[7:0];
  _RAND_6009 = {1{`RANDOM}};
  lineBuffer_6002 = _RAND_6009[7:0];
  _RAND_6010 = {1{`RANDOM}};
  lineBuffer_6003 = _RAND_6010[7:0];
  _RAND_6011 = {1{`RANDOM}};
  lineBuffer_6004 = _RAND_6011[7:0];
  _RAND_6012 = {1{`RANDOM}};
  lineBuffer_6005 = _RAND_6012[7:0];
  _RAND_6013 = {1{`RANDOM}};
  lineBuffer_6006 = _RAND_6013[7:0];
  _RAND_6014 = {1{`RANDOM}};
  lineBuffer_6007 = _RAND_6014[7:0];
  _RAND_6015 = {1{`RANDOM}};
  lineBuffer_6008 = _RAND_6015[7:0];
  _RAND_6016 = {1{`RANDOM}};
  lineBuffer_6009 = _RAND_6016[7:0];
  _RAND_6017 = {1{`RANDOM}};
  lineBuffer_6010 = _RAND_6017[7:0];
  _RAND_6018 = {1{`RANDOM}};
  lineBuffer_6011 = _RAND_6018[7:0];
  _RAND_6019 = {1{`RANDOM}};
  lineBuffer_6012 = _RAND_6019[7:0];
  _RAND_6020 = {1{`RANDOM}};
  lineBuffer_6013 = _RAND_6020[7:0];
  _RAND_6021 = {1{`RANDOM}};
  lineBuffer_6014 = _RAND_6021[7:0];
  _RAND_6022 = {1{`RANDOM}};
  lineBuffer_6015 = _RAND_6022[7:0];
  _RAND_6023 = {1{`RANDOM}};
  lineBuffer_6016 = _RAND_6023[7:0];
  _RAND_6024 = {1{`RANDOM}};
  lineBuffer_6017 = _RAND_6024[7:0];
  _RAND_6025 = {1{`RANDOM}};
  lineBuffer_6018 = _RAND_6025[7:0];
  _RAND_6026 = {1{`RANDOM}};
  lineBuffer_6019 = _RAND_6026[7:0];
  _RAND_6027 = {1{`RANDOM}};
  lineBuffer_6020 = _RAND_6027[7:0];
  _RAND_6028 = {1{`RANDOM}};
  lineBuffer_6021 = _RAND_6028[7:0];
  _RAND_6029 = {1{`RANDOM}};
  lineBuffer_6022 = _RAND_6029[7:0];
  _RAND_6030 = {1{`RANDOM}};
  lineBuffer_6023 = _RAND_6030[7:0];
  _RAND_6031 = {1{`RANDOM}};
  lineBuffer_6024 = _RAND_6031[7:0];
  _RAND_6032 = {1{`RANDOM}};
  lineBuffer_6025 = _RAND_6032[7:0];
  _RAND_6033 = {1{`RANDOM}};
  lineBuffer_6026 = _RAND_6033[7:0];
  _RAND_6034 = {1{`RANDOM}};
  lineBuffer_6027 = _RAND_6034[7:0];
  _RAND_6035 = {1{`RANDOM}};
  lineBuffer_6028 = _RAND_6035[7:0];
  _RAND_6036 = {1{`RANDOM}};
  lineBuffer_6029 = _RAND_6036[7:0];
  _RAND_6037 = {1{`RANDOM}};
  lineBuffer_6030 = _RAND_6037[7:0];
  _RAND_6038 = {1{`RANDOM}};
  lineBuffer_6031 = _RAND_6038[7:0];
  _RAND_6039 = {1{`RANDOM}};
  lineBuffer_6032 = _RAND_6039[7:0];
  _RAND_6040 = {1{`RANDOM}};
  lineBuffer_6033 = _RAND_6040[7:0];
  _RAND_6041 = {1{`RANDOM}};
  lineBuffer_6034 = _RAND_6041[7:0];
  _RAND_6042 = {1{`RANDOM}};
  lineBuffer_6035 = _RAND_6042[7:0];
  _RAND_6043 = {1{`RANDOM}};
  lineBuffer_6036 = _RAND_6043[7:0];
  _RAND_6044 = {1{`RANDOM}};
  lineBuffer_6037 = _RAND_6044[7:0];
  _RAND_6045 = {1{`RANDOM}};
  lineBuffer_6038 = _RAND_6045[7:0];
  _RAND_6046 = {1{`RANDOM}};
  lineBuffer_6039 = _RAND_6046[7:0];
  _RAND_6047 = {1{`RANDOM}};
  lineBuffer_6040 = _RAND_6047[7:0];
  _RAND_6048 = {1{`RANDOM}};
  lineBuffer_6041 = _RAND_6048[7:0];
  _RAND_6049 = {1{`RANDOM}};
  lineBuffer_6042 = _RAND_6049[7:0];
  _RAND_6050 = {1{`RANDOM}};
  lineBuffer_6043 = _RAND_6050[7:0];
  _RAND_6051 = {1{`RANDOM}};
  lineBuffer_6044 = _RAND_6051[7:0];
  _RAND_6052 = {1{`RANDOM}};
  lineBuffer_6045 = _RAND_6052[7:0];
  _RAND_6053 = {1{`RANDOM}};
  lineBuffer_6046 = _RAND_6053[7:0];
  _RAND_6054 = {1{`RANDOM}};
  lineBuffer_6047 = _RAND_6054[7:0];
  _RAND_6055 = {1{`RANDOM}};
  lineBuffer_6048 = _RAND_6055[7:0];
  _RAND_6056 = {1{`RANDOM}};
  lineBuffer_6049 = _RAND_6056[7:0];
  _RAND_6057 = {1{`RANDOM}};
  lineBuffer_6050 = _RAND_6057[7:0];
  _RAND_6058 = {1{`RANDOM}};
  lineBuffer_6051 = _RAND_6058[7:0];
  _RAND_6059 = {1{`RANDOM}};
  lineBuffer_6052 = _RAND_6059[7:0];
  _RAND_6060 = {1{`RANDOM}};
  lineBuffer_6053 = _RAND_6060[7:0];
  _RAND_6061 = {1{`RANDOM}};
  lineBuffer_6054 = _RAND_6061[7:0];
  _RAND_6062 = {1{`RANDOM}};
  lineBuffer_6055 = _RAND_6062[7:0];
  _RAND_6063 = {1{`RANDOM}};
  lineBuffer_6056 = _RAND_6063[7:0];
  _RAND_6064 = {1{`RANDOM}};
  lineBuffer_6057 = _RAND_6064[7:0];
  _RAND_6065 = {1{`RANDOM}};
  lineBuffer_6058 = _RAND_6065[7:0];
  _RAND_6066 = {1{`RANDOM}};
  lineBuffer_6059 = _RAND_6066[7:0];
  _RAND_6067 = {1{`RANDOM}};
  lineBuffer_6060 = _RAND_6067[7:0];
  _RAND_6068 = {1{`RANDOM}};
  lineBuffer_6061 = _RAND_6068[7:0];
  _RAND_6069 = {1{`RANDOM}};
  lineBuffer_6062 = _RAND_6069[7:0];
  _RAND_6070 = {1{`RANDOM}};
  lineBuffer_6063 = _RAND_6070[7:0];
  _RAND_6071 = {1{`RANDOM}};
  lineBuffer_6064 = _RAND_6071[7:0];
  _RAND_6072 = {1{`RANDOM}};
  lineBuffer_6065 = _RAND_6072[7:0];
  _RAND_6073 = {1{`RANDOM}};
  lineBuffer_6066 = _RAND_6073[7:0];
  _RAND_6074 = {1{`RANDOM}};
  lineBuffer_6067 = _RAND_6074[7:0];
  _RAND_6075 = {1{`RANDOM}};
  lineBuffer_6068 = _RAND_6075[7:0];
  _RAND_6076 = {1{`RANDOM}};
  lineBuffer_6069 = _RAND_6076[7:0];
  _RAND_6077 = {1{`RANDOM}};
  lineBuffer_6070 = _RAND_6077[7:0];
  _RAND_6078 = {1{`RANDOM}};
  lineBuffer_6071 = _RAND_6078[7:0];
  _RAND_6079 = {1{`RANDOM}};
  lineBuffer_6072 = _RAND_6079[7:0];
  _RAND_6080 = {1{`RANDOM}};
  lineBuffer_6073 = _RAND_6080[7:0];
  _RAND_6081 = {1{`RANDOM}};
  lineBuffer_6074 = _RAND_6081[7:0];
  _RAND_6082 = {1{`RANDOM}};
  lineBuffer_6075 = _RAND_6082[7:0];
  _RAND_6083 = {1{`RANDOM}};
  lineBuffer_6076 = _RAND_6083[7:0];
  _RAND_6084 = {1{`RANDOM}};
  lineBuffer_6077 = _RAND_6084[7:0];
  _RAND_6085 = {1{`RANDOM}};
  lineBuffer_6078 = _RAND_6085[7:0];
  _RAND_6086 = {1{`RANDOM}};
  lineBuffer_6079 = _RAND_6086[7:0];
  _RAND_6087 = {1{`RANDOM}};
  lineBuffer_6080 = _RAND_6087[7:0];
  _RAND_6088 = {1{`RANDOM}};
  lineBuffer_6081 = _RAND_6088[7:0];
  _RAND_6089 = {1{`RANDOM}};
  lineBuffer_6082 = _RAND_6089[7:0];
  _RAND_6090 = {1{`RANDOM}};
  lineBuffer_6083 = _RAND_6090[7:0];
  _RAND_6091 = {1{`RANDOM}};
  lineBuffer_6084 = _RAND_6091[7:0];
  _RAND_6092 = {1{`RANDOM}};
  lineBuffer_6085 = _RAND_6092[7:0];
  _RAND_6093 = {1{`RANDOM}};
  lineBuffer_6086 = _RAND_6093[7:0];
  _RAND_6094 = {1{`RANDOM}};
  lineBuffer_6087 = _RAND_6094[7:0];
  _RAND_6095 = {1{`RANDOM}};
  lineBuffer_6088 = _RAND_6095[7:0];
  _RAND_6096 = {1{`RANDOM}};
  lineBuffer_6089 = _RAND_6096[7:0];
  _RAND_6097 = {1{`RANDOM}};
  lineBuffer_6090 = _RAND_6097[7:0];
  _RAND_6098 = {1{`RANDOM}};
  lineBuffer_6091 = _RAND_6098[7:0];
  _RAND_6099 = {1{`RANDOM}};
  lineBuffer_6092 = _RAND_6099[7:0];
  _RAND_6100 = {1{`RANDOM}};
  lineBuffer_6093 = _RAND_6100[7:0];
  _RAND_6101 = {1{`RANDOM}};
  lineBuffer_6094 = _RAND_6101[7:0];
  _RAND_6102 = {1{`RANDOM}};
  lineBuffer_6095 = _RAND_6102[7:0];
  _RAND_6103 = {1{`RANDOM}};
  lineBuffer_6096 = _RAND_6103[7:0];
  _RAND_6104 = {1{`RANDOM}};
  lineBuffer_6097 = _RAND_6104[7:0];
  _RAND_6105 = {1{`RANDOM}};
  lineBuffer_6098 = _RAND_6105[7:0];
  _RAND_6106 = {1{`RANDOM}};
  lineBuffer_6099 = _RAND_6106[7:0];
  _RAND_6107 = {1{`RANDOM}};
  lineBuffer_6100 = _RAND_6107[7:0];
  _RAND_6108 = {1{`RANDOM}};
  lineBuffer_6101 = _RAND_6108[7:0];
  _RAND_6109 = {1{`RANDOM}};
  lineBuffer_6102 = _RAND_6109[7:0];
  _RAND_6110 = {1{`RANDOM}};
  lineBuffer_6103 = _RAND_6110[7:0];
  _RAND_6111 = {1{`RANDOM}};
  lineBuffer_6104 = _RAND_6111[7:0];
  _RAND_6112 = {1{`RANDOM}};
  lineBuffer_6105 = _RAND_6112[7:0];
  _RAND_6113 = {1{`RANDOM}};
  lineBuffer_6106 = _RAND_6113[7:0];
  _RAND_6114 = {1{`RANDOM}};
  lineBuffer_6107 = _RAND_6114[7:0];
  _RAND_6115 = {1{`RANDOM}};
  lineBuffer_6108 = _RAND_6115[7:0];
  _RAND_6116 = {1{`RANDOM}};
  lineBuffer_6109 = _RAND_6116[7:0];
  _RAND_6117 = {1{`RANDOM}};
  lineBuffer_6110 = _RAND_6117[7:0];
  _RAND_6118 = {1{`RANDOM}};
  lineBuffer_6111 = _RAND_6118[7:0];
  _RAND_6119 = {1{`RANDOM}};
  lineBuffer_6112 = _RAND_6119[7:0];
  _RAND_6120 = {1{`RANDOM}};
  lineBuffer_6113 = _RAND_6120[7:0];
  _RAND_6121 = {1{`RANDOM}};
  lineBuffer_6114 = _RAND_6121[7:0];
  _RAND_6122 = {1{`RANDOM}};
  lineBuffer_6115 = _RAND_6122[7:0];
  _RAND_6123 = {1{`RANDOM}};
  lineBuffer_6116 = _RAND_6123[7:0];
  _RAND_6124 = {1{`RANDOM}};
  lineBuffer_6117 = _RAND_6124[7:0];
  _RAND_6125 = {1{`RANDOM}};
  lineBuffer_6118 = _RAND_6125[7:0];
  _RAND_6126 = {1{`RANDOM}};
  lineBuffer_6119 = _RAND_6126[7:0];
  _RAND_6127 = {1{`RANDOM}};
  lineBuffer_6120 = _RAND_6127[7:0];
  _RAND_6128 = {1{`RANDOM}};
  lineBuffer_6121 = _RAND_6128[7:0];
  _RAND_6129 = {1{`RANDOM}};
  lineBuffer_6122 = _RAND_6129[7:0];
  _RAND_6130 = {1{`RANDOM}};
  lineBuffer_6123 = _RAND_6130[7:0];
  _RAND_6131 = {1{`RANDOM}};
  lineBuffer_6124 = _RAND_6131[7:0];
  _RAND_6132 = {1{`RANDOM}};
  lineBuffer_6125 = _RAND_6132[7:0];
  _RAND_6133 = {1{`RANDOM}};
  lineBuffer_6126 = _RAND_6133[7:0];
  _RAND_6134 = {1{`RANDOM}};
  lineBuffer_6127 = _RAND_6134[7:0];
  _RAND_6135 = {1{`RANDOM}};
  lineBuffer_6128 = _RAND_6135[7:0];
  _RAND_6136 = {1{`RANDOM}};
  lineBuffer_6129 = _RAND_6136[7:0];
  _RAND_6137 = {1{`RANDOM}};
  lineBuffer_6130 = _RAND_6137[7:0];
  _RAND_6138 = {1{`RANDOM}};
  lineBuffer_6131 = _RAND_6138[7:0];
  _RAND_6139 = {1{`RANDOM}};
  lineBuffer_6132 = _RAND_6139[7:0];
  _RAND_6140 = {1{`RANDOM}};
  lineBuffer_6133 = _RAND_6140[7:0];
  _RAND_6141 = {1{`RANDOM}};
  lineBuffer_6134 = _RAND_6141[7:0];
  _RAND_6142 = {1{`RANDOM}};
  lineBuffer_6135 = _RAND_6142[7:0];
  _RAND_6143 = {1{`RANDOM}};
  lineBuffer_6136 = _RAND_6143[7:0];
  _RAND_6144 = {1{`RANDOM}};
  lineBuffer_6137 = _RAND_6144[7:0];
  _RAND_6145 = {1{`RANDOM}};
  lineBuffer_6138 = _RAND_6145[7:0];
  _RAND_6146 = {1{`RANDOM}};
  lineBuffer_6139 = _RAND_6146[7:0];
  _RAND_6147 = {1{`RANDOM}};
  lineBuffer_6140 = _RAND_6147[7:0];
  _RAND_6148 = {1{`RANDOM}};
  lineBuffer_6141 = _RAND_6148[7:0];
  _RAND_6149 = {1{`RANDOM}};
  lineBuffer_6142 = _RAND_6149[7:0];
  _RAND_6150 = {1{`RANDOM}};
  lineBuffer_6143 = _RAND_6150[7:0];
  _RAND_6151 = {1{`RANDOM}};
  lineBuffer_6144 = _RAND_6151[7:0];
  _RAND_6152 = {1{`RANDOM}};
  lineBuffer_6145 = _RAND_6152[7:0];
  _RAND_6153 = {1{`RANDOM}};
  lineBuffer_6146 = _RAND_6153[7:0];
  _RAND_6154 = {1{`RANDOM}};
  lineBuffer_6147 = _RAND_6154[7:0];
  _RAND_6155 = {1{`RANDOM}};
  lineBuffer_6148 = _RAND_6155[7:0];
  _RAND_6156 = {1{`RANDOM}};
  lineBuffer_6149 = _RAND_6156[7:0];
  _RAND_6157 = {1{`RANDOM}};
  lineBuffer_6150 = _RAND_6157[7:0];
  _RAND_6158 = {1{`RANDOM}};
  lineBuffer_6151 = _RAND_6158[7:0];
  _RAND_6159 = {1{`RANDOM}};
  lineBuffer_6152 = _RAND_6159[7:0];
  _RAND_6160 = {1{`RANDOM}};
  lineBuffer_6153 = _RAND_6160[7:0];
  _RAND_6161 = {1{`RANDOM}};
  lineBuffer_6154 = _RAND_6161[7:0];
  _RAND_6162 = {1{`RANDOM}};
  lineBuffer_6155 = _RAND_6162[7:0];
  _RAND_6163 = {1{`RANDOM}};
  lineBuffer_6156 = _RAND_6163[7:0];
  _RAND_6164 = {1{`RANDOM}};
  lineBuffer_6157 = _RAND_6164[7:0];
  _RAND_6165 = {1{`RANDOM}};
  lineBuffer_6158 = _RAND_6165[7:0];
  _RAND_6166 = {1{`RANDOM}};
  lineBuffer_6159 = _RAND_6166[7:0];
  _RAND_6167 = {1{`RANDOM}};
  lineBuffer_6160 = _RAND_6167[7:0];
  _RAND_6168 = {1{`RANDOM}};
  lineBuffer_6161 = _RAND_6168[7:0];
  _RAND_6169 = {1{`RANDOM}};
  lineBuffer_6162 = _RAND_6169[7:0];
  _RAND_6170 = {1{`RANDOM}};
  lineBuffer_6163 = _RAND_6170[7:0];
  _RAND_6171 = {1{`RANDOM}};
  lineBuffer_6164 = _RAND_6171[7:0];
  _RAND_6172 = {1{`RANDOM}};
  lineBuffer_6165 = _RAND_6172[7:0];
  _RAND_6173 = {1{`RANDOM}};
  lineBuffer_6166 = _RAND_6173[7:0];
  _RAND_6174 = {1{`RANDOM}};
  lineBuffer_6167 = _RAND_6174[7:0];
  _RAND_6175 = {1{`RANDOM}};
  lineBuffer_6168 = _RAND_6175[7:0];
  _RAND_6176 = {1{`RANDOM}};
  lineBuffer_6169 = _RAND_6176[7:0];
  _RAND_6177 = {1{`RANDOM}};
  lineBuffer_6170 = _RAND_6177[7:0];
  _RAND_6178 = {1{`RANDOM}};
  lineBuffer_6171 = _RAND_6178[7:0];
  _RAND_6179 = {1{`RANDOM}};
  lineBuffer_6172 = _RAND_6179[7:0];
  _RAND_6180 = {1{`RANDOM}};
  lineBuffer_6173 = _RAND_6180[7:0];
  _RAND_6181 = {1{`RANDOM}};
  lineBuffer_6174 = _RAND_6181[7:0];
  _RAND_6182 = {1{`RANDOM}};
  lineBuffer_6175 = _RAND_6182[7:0];
  _RAND_6183 = {1{`RANDOM}};
  lineBuffer_6176 = _RAND_6183[7:0];
  _RAND_6184 = {1{`RANDOM}};
  lineBuffer_6177 = _RAND_6184[7:0];
  _RAND_6185 = {1{`RANDOM}};
  lineBuffer_6178 = _RAND_6185[7:0];
  _RAND_6186 = {1{`RANDOM}};
  lineBuffer_6179 = _RAND_6186[7:0];
  _RAND_6187 = {1{`RANDOM}};
  lineBuffer_6180 = _RAND_6187[7:0];
  _RAND_6188 = {1{`RANDOM}};
  lineBuffer_6181 = _RAND_6188[7:0];
  _RAND_6189 = {1{`RANDOM}};
  lineBuffer_6182 = _RAND_6189[7:0];
  _RAND_6190 = {1{`RANDOM}};
  lineBuffer_6183 = _RAND_6190[7:0];
  _RAND_6191 = {1{`RANDOM}};
  lineBuffer_6184 = _RAND_6191[7:0];
  _RAND_6192 = {1{`RANDOM}};
  lineBuffer_6185 = _RAND_6192[7:0];
  _RAND_6193 = {1{`RANDOM}};
  lineBuffer_6186 = _RAND_6193[7:0];
  _RAND_6194 = {1{`RANDOM}};
  lineBuffer_6187 = _RAND_6194[7:0];
  _RAND_6195 = {1{`RANDOM}};
  lineBuffer_6188 = _RAND_6195[7:0];
  _RAND_6196 = {1{`RANDOM}};
  lineBuffer_6189 = _RAND_6196[7:0];
  _RAND_6197 = {1{`RANDOM}};
  lineBuffer_6190 = _RAND_6197[7:0];
  _RAND_6198 = {1{`RANDOM}};
  lineBuffer_6191 = _RAND_6198[7:0];
  _RAND_6199 = {1{`RANDOM}};
  lineBuffer_6192 = _RAND_6199[7:0];
  _RAND_6200 = {1{`RANDOM}};
  lineBuffer_6193 = _RAND_6200[7:0];
  _RAND_6201 = {1{`RANDOM}};
  lineBuffer_6194 = _RAND_6201[7:0];
  _RAND_6202 = {1{`RANDOM}};
  lineBuffer_6195 = _RAND_6202[7:0];
  _RAND_6203 = {1{`RANDOM}};
  lineBuffer_6196 = _RAND_6203[7:0];
  _RAND_6204 = {1{`RANDOM}};
  lineBuffer_6197 = _RAND_6204[7:0];
  _RAND_6205 = {1{`RANDOM}};
  lineBuffer_6198 = _RAND_6205[7:0];
  _RAND_6206 = {1{`RANDOM}};
  lineBuffer_6199 = _RAND_6206[7:0];
  _RAND_6207 = {1{`RANDOM}};
  lineBuffer_6200 = _RAND_6207[7:0];
  _RAND_6208 = {1{`RANDOM}};
  lineBuffer_6201 = _RAND_6208[7:0];
  _RAND_6209 = {1{`RANDOM}};
  lineBuffer_6202 = _RAND_6209[7:0];
  _RAND_6210 = {1{`RANDOM}};
  lineBuffer_6203 = _RAND_6210[7:0];
  _RAND_6211 = {1{`RANDOM}};
  lineBuffer_6204 = _RAND_6211[7:0];
  _RAND_6212 = {1{`RANDOM}};
  lineBuffer_6205 = _RAND_6212[7:0];
  _RAND_6213 = {1{`RANDOM}};
  lineBuffer_6206 = _RAND_6213[7:0];
  _RAND_6214 = {1{`RANDOM}};
  lineBuffer_6207 = _RAND_6214[7:0];
  _RAND_6215 = {1{`RANDOM}};
  lineBuffer_6208 = _RAND_6215[7:0];
  _RAND_6216 = {1{`RANDOM}};
  lineBuffer_6209 = _RAND_6216[7:0];
  _RAND_6217 = {1{`RANDOM}};
  lineBuffer_6210 = _RAND_6217[7:0];
  _RAND_6218 = {1{`RANDOM}};
  lineBuffer_6211 = _RAND_6218[7:0];
  _RAND_6219 = {1{`RANDOM}};
  lineBuffer_6212 = _RAND_6219[7:0];
  _RAND_6220 = {1{`RANDOM}};
  lineBuffer_6213 = _RAND_6220[7:0];
  _RAND_6221 = {1{`RANDOM}};
  lineBuffer_6214 = _RAND_6221[7:0];
  _RAND_6222 = {1{`RANDOM}};
  lineBuffer_6215 = _RAND_6222[7:0];
  _RAND_6223 = {1{`RANDOM}};
  lineBuffer_6216 = _RAND_6223[7:0];
  _RAND_6224 = {1{`RANDOM}};
  lineBuffer_6217 = _RAND_6224[7:0];
  _RAND_6225 = {1{`RANDOM}};
  lineBuffer_6218 = _RAND_6225[7:0];
  _RAND_6226 = {1{`RANDOM}};
  lineBuffer_6219 = _RAND_6226[7:0];
  _RAND_6227 = {1{`RANDOM}};
  lineBuffer_6220 = _RAND_6227[7:0];
  _RAND_6228 = {1{`RANDOM}};
  lineBuffer_6221 = _RAND_6228[7:0];
  _RAND_6229 = {1{`RANDOM}};
  lineBuffer_6222 = _RAND_6229[7:0];
  _RAND_6230 = {1{`RANDOM}};
  lineBuffer_6223 = _RAND_6230[7:0];
  _RAND_6231 = {1{`RANDOM}};
  lineBuffer_6224 = _RAND_6231[7:0];
  _RAND_6232 = {1{`RANDOM}};
  lineBuffer_6225 = _RAND_6232[7:0];
  _RAND_6233 = {1{`RANDOM}};
  lineBuffer_6226 = _RAND_6233[7:0];
  _RAND_6234 = {1{`RANDOM}};
  lineBuffer_6227 = _RAND_6234[7:0];
  _RAND_6235 = {1{`RANDOM}};
  lineBuffer_6228 = _RAND_6235[7:0];
  _RAND_6236 = {1{`RANDOM}};
  lineBuffer_6229 = _RAND_6236[7:0];
  _RAND_6237 = {1{`RANDOM}};
  lineBuffer_6230 = _RAND_6237[7:0];
  _RAND_6238 = {1{`RANDOM}};
  lineBuffer_6231 = _RAND_6238[7:0];
  _RAND_6239 = {1{`RANDOM}};
  lineBuffer_6232 = _RAND_6239[7:0];
  _RAND_6240 = {1{`RANDOM}};
  lineBuffer_6233 = _RAND_6240[7:0];
  _RAND_6241 = {1{`RANDOM}};
  lineBuffer_6234 = _RAND_6241[7:0];
  _RAND_6242 = {1{`RANDOM}};
  lineBuffer_6235 = _RAND_6242[7:0];
  _RAND_6243 = {1{`RANDOM}};
  lineBuffer_6236 = _RAND_6243[7:0];
  _RAND_6244 = {1{`RANDOM}};
  lineBuffer_6237 = _RAND_6244[7:0];
  _RAND_6245 = {1{`RANDOM}};
  lineBuffer_6238 = _RAND_6245[7:0];
  _RAND_6246 = {1{`RANDOM}};
  lineBuffer_6239 = _RAND_6246[7:0];
  _RAND_6247 = {1{`RANDOM}};
  lineBuffer_6240 = _RAND_6247[7:0];
  _RAND_6248 = {1{`RANDOM}};
  lineBuffer_6241 = _RAND_6248[7:0];
  _RAND_6249 = {1{`RANDOM}};
  lineBuffer_6242 = _RAND_6249[7:0];
  _RAND_6250 = {1{`RANDOM}};
  lineBuffer_6243 = _RAND_6250[7:0];
  _RAND_6251 = {1{`RANDOM}};
  lineBuffer_6244 = _RAND_6251[7:0];
  _RAND_6252 = {1{`RANDOM}};
  lineBuffer_6245 = _RAND_6252[7:0];
  _RAND_6253 = {1{`RANDOM}};
  lineBuffer_6246 = _RAND_6253[7:0];
  _RAND_6254 = {1{`RANDOM}};
  lineBuffer_6247 = _RAND_6254[7:0];
  _RAND_6255 = {1{`RANDOM}};
  lineBuffer_6248 = _RAND_6255[7:0];
  _RAND_6256 = {1{`RANDOM}};
  lineBuffer_6249 = _RAND_6256[7:0];
  _RAND_6257 = {1{`RANDOM}};
  lineBuffer_6250 = _RAND_6257[7:0];
  _RAND_6258 = {1{`RANDOM}};
  lineBuffer_6251 = _RAND_6258[7:0];
  _RAND_6259 = {1{`RANDOM}};
  lineBuffer_6252 = _RAND_6259[7:0];
  _RAND_6260 = {1{`RANDOM}};
  lineBuffer_6253 = _RAND_6260[7:0];
  _RAND_6261 = {1{`RANDOM}};
  lineBuffer_6254 = _RAND_6261[7:0];
  _RAND_6262 = {1{`RANDOM}};
  lineBuffer_6255 = _RAND_6262[7:0];
  _RAND_6263 = {1{`RANDOM}};
  lineBuffer_6256 = _RAND_6263[7:0];
  _RAND_6264 = {1{`RANDOM}};
  lineBuffer_6257 = _RAND_6264[7:0];
  _RAND_6265 = {1{`RANDOM}};
  lineBuffer_6258 = _RAND_6265[7:0];
  _RAND_6266 = {1{`RANDOM}};
  lineBuffer_6259 = _RAND_6266[7:0];
  _RAND_6267 = {1{`RANDOM}};
  lineBuffer_6260 = _RAND_6267[7:0];
  _RAND_6268 = {1{`RANDOM}};
  lineBuffer_6261 = _RAND_6268[7:0];
  _RAND_6269 = {1{`RANDOM}};
  lineBuffer_6262 = _RAND_6269[7:0];
  _RAND_6270 = {1{`RANDOM}};
  lineBuffer_6263 = _RAND_6270[7:0];
  _RAND_6271 = {1{`RANDOM}};
  lineBuffer_6264 = _RAND_6271[7:0];
  _RAND_6272 = {1{`RANDOM}};
  lineBuffer_6265 = _RAND_6272[7:0];
  _RAND_6273 = {1{`RANDOM}};
  lineBuffer_6266 = _RAND_6273[7:0];
  _RAND_6274 = {1{`RANDOM}};
  lineBuffer_6267 = _RAND_6274[7:0];
  _RAND_6275 = {1{`RANDOM}};
  lineBuffer_6268 = _RAND_6275[7:0];
  _RAND_6276 = {1{`RANDOM}};
  lineBuffer_6269 = _RAND_6276[7:0];
  _RAND_6277 = {1{`RANDOM}};
  lineBuffer_6270 = _RAND_6277[7:0];
  _RAND_6278 = {1{`RANDOM}};
  lineBuffer_6271 = _RAND_6278[7:0];
  _RAND_6279 = {1{`RANDOM}};
  lineBuffer_6272 = _RAND_6279[7:0];
  _RAND_6280 = {1{`RANDOM}};
  lineBuffer_6273 = _RAND_6280[7:0];
  _RAND_6281 = {1{`RANDOM}};
  lineBuffer_6274 = _RAND_6281[7:0];
  _RAND_6282 = {1{`RANDOM}};
  lineBuffer_6275 = _RAND_6282[7:0];
  _RAND_6283 = {1{`RANDOM}};
  lineBuffer_6276 = _RAND_6283[7:0];
  _RAND_6284 = {1{`RANDOM}};
  lineBuffer_6277 = _RAND_6284[7:0];
  _RAND_6285 = {1{`RANDOM}};
  lineBuffer_6278 = _RAND_6285[7:0];
  _RAND_6286 = {1{`RANDOM}};
  lineBuffer_6279 = _RAND_6286[7:0];
  _RAND_6287 = {1{`RANDOM}};
  lineBuffer_6280 = _RAND_6287[7:0];
  _RAND_6288 = {1{`RANDOM}};
  lineBuffer_6281 = _RAND_6288[7:0];
  _RAND_6289 = {1{`RANDOM}};
  lineBuffer_6282 = _RAND_6289[7:0];
  _RAND_6290 = {1{`RANDOM}};
  lineBuffer_6283 = _RAND_6290[7:0];
  _RAND_6291 = {1{`RANDOM}};
  lineBuffer_6284 = _RAND_6291[7:0];
  _RAND_6292 = {1{`RANDOM}};
  lineBuffer_6285 = _RAND_6292[7:0];
  _RAND_6293 = {1{`RANDOM}};
  lineBuffer_6286 = _RAND_6293[7:0];
  _RAND_6294 = {1{`RANDOM}};
  lineBuffer_6287 = _RAND_6294[7:0];
  _RAND_6295 = {1{`RANDOM}};
  lineBuffer_6288 = _RAND_6295[7:0];
  _RAND_6296 = {1{`RANDOM}};
  lineBuffer_6289 = _RAND_6296[7:0];
  _RAND_6297 = {1{`RANDOM}};
  lineBuffer_6290 = _RAND_6297[7:0];
  _RAND_6298 = {1{`RANDOM}};
  lineBuffer_6291 = _RAND_6298[7:0];
  _RAND_6299 = {1{`RANDOM}};
  lineBuffer_6292 = _RAND_6299[7:0];
  _RAND_6300 = {1{`RANDOM}};
  lineBuffer_6293 = _RAND_6300[7:0];
  _RAND_6301 = {1{`RANDOM}};
  lineBuffer_6294 = _RAND_6301[7:0];
  _RAND_6302 = {1{`RANDOM}};
  lineBuffer_6295 = _RAND_6302[7:0];
  _RAND_6303 = {1{`RANDOM}};
  lineBuffer_6296 = _RAND_6303[7:0];
  _RAND_6304 = {1{`RANDOM}};
  lineBuffer_6297 = _RAND_6304[7:0];
  _RAND_6305 = {1{`RANDOM}};
  lineBuffer_6298 = _RAND_6305[7:0];
  _RAND_6306 = {1{`RANDOM}};
  lineBuffer_6299 = _RAND_6306[7:0];
  _RAND_6307 = {1{`RANDOM}};
  lineBuffer_6300 = _RAND_6307[7:0];
  _RAND_6308 = {1{`RANDOM}};
  lineBuffer_6301 = _RAND_6308[7:0];
  _RAND_6309 = {1{`RANDOM}};
  lineBuffer_6302 = _RAND_6309[7:0];
  _RAND_6310 = {1{`RANDOM}};
  lineBuffer_6303 = _RAND_6310[7:0];
  _RAND_6311 = {1{`RANDOM}};
  lineBuffer_6304 = _RAND_6311[7:0];
  _RAND_6312 = {1{`RANDOM}};
  lineBuffer_6305 = _RAND_6312[7:0];
  _RAND_6313 = {1{`RANDOM}};
  lineBuffer_6306 = _RAND_6313[7:0];
  _RAND_6314 = {1{`RANDOM}};
  lineBuffer_6307 = _RAND_6314[7:0];
  _RAND_6315 = {1{`RANDOM}};
  lineBuffer_6308 = _RAND_6315[7:0];
  _RAND_6316 = {1{`RANDOM}};
  lineBuffer_6309 = _RAND_6316[7:0];
  _RAND_6317 = {1{`RANDOM}};
  lineBuffer_6310 = _RAND_6317[7:0];
  _RAND_6318 = {1{`RANDOM}};
  lineBuffer_6311 = _RAND_6318[7:0];
  _RAND_6319 = {1{`RANDOM}};
  lineBuffer_6312 = _RAND_6319[7:0];
  _RAND_6320 = {1{`RANDOM}};
  lineBuffer_6313 = _RAND_6320[7:0];
  _RAND_6321 = {1{`RANDOM}};
  lineBuffer_6314 = _RAND_6321[7:0];
  _RAND_6322 = {1{`RANDOM}};
  lineBuffer_6315 = _RAND_6322[7:0];
  _RAND_6323 = {1{`RANDOM}};
  lineBuffer_6316 = _RAND_6323[7:0];
  _RAND_6324 = {1{`RANDOM}};
  lineBuffer_6317 = _RAND_6324[7:0];
  _RAND_6325 = {1{`RANDOM}};
  lineBuffer_6318 = _RAND_6325[7:0];
  _RAND_6326 = {1{`RANDOM}};
  lineBuffer_6319 = _RAND_6326[7:0];
  _RAND_6327 = {1{`RANDOM}};
  lineBuffer_6320 = _RAND_6327[7:0];
  _RAND_6328 = {1{`RANDOM}};
  lineBuffer_6321 = _RAND_6328[7:0];
  _RAND_6329 = {1{`RANDOM}};
  lineBuffer_6322 = _RAND_6329[7:0];
  _RAND_6330 = {1{`RANDOM}};
  lineBuffer_6323 = _RAND_6330[7:0];
  _RAND_6331 = {1{`RANDOM}};
  lineBuffer_6324 = _RAND_6331[7:0];
  _RAND_6332 = {1{`RANDOM}};
  lineBuffer_6325 = _RAND_6332[7:0];
  _RAND_6333 = {1{`RANDOM}};
  lineBuffer_6326 = _RAND_6333[7:0];
  _RAND_6334 = {1{`RANDOM}};
  lineBuffer_6327 = _RAND_6334[7:0];
  _RAND_6335 = {1{`RANDOM}};
  lineBuffer_6328 = _RAND_6335[7:0];
  _RAND_6336 = {1{`RANDOM}};
  lineBuffer_6329 = _RAND_6336[7:0];
  _RAND_6337 = {1{`RANDOM}};
  lineBuffer_6330 = _RAND_6337[7:0];
  _RAND_6338 = {1{`RANDOM}};
  lineBuffer_6331 = _RAND_6338[7:0];
  _RAND_6339 = {1{`RANDOM}};
  lineBuffer_6332 = _RAND_6339[7:0];
  _RAND_6340 = {1{`RANDOM}};
  lineBuffer_6333 = _RAND_6340[7:0];
  _RAND_6341 = {1{`RANDOM}};
  lineBuffer_6334 = _RAND_6341[7:0];
  _RAND_6342 = {1{`RANDOM}};
  lineBuffer_6335 = _RAND_6342[7:0];
  _RAND_6343 = {1{`RANDOM}};
  lineBuffer_6336 = _RAND_6343[7:0];
  _RAND_6344 = {1{`RANDOM}};
  lineBuffer_6337 = _RAND_6344[7:0];
  _RAND_6345 = {1{`RANDOM}};
  lineBuffer_6338 = _RAND_6345[7:0];
  _RAND_6346 = {1{`RANDOM}};
  lineBuffer_6339 = _RAND_6346[7:0];
  _RAND_6347 = {1{`RANDOM}};
  lineBuffer_6340 = _RAND_6347[7:0];
  _RAND_6348 = {1{`RANDOM}};
  lineBuffer_6341 = _RAND_6348[7:0];
  _RAND_6349 = {1{`RANDOM}};
  lineBuffer_6342 = _RAND_6349[7:0];
  _RAND_6350 = {1{`RANDOM}};
  lineBuffer_6343 = _RAND_6350[7:0];
  _RAND_6351 = {1{`RANDOM}};
  lineBuffer_6344 = _RAND_6351[7:0];
  _RAND_6352 = {1{`RANDOM}};
  lineBuffer_6345 = _RAND_6352[7:0];
  _RAND_6353 = {1{`RANDOM}};
  lineBuffer_6346 = _RAND_6353[7:0];
  _RAND_6354 = {1{`RANDOM}};
  lineBuffer_6347 = _RAND_6354[7:0];
  _RAND_6355 = {1{`RANDOM}};
  lineBuffer_6348 = _RAND_6355[7:0];
  _RAND_6356 = {1{`RANDOM}};
  lineBuffer_6349 = _RAND_6356[7:0];
  _RAND_6357 = {1{`RANDOM}};
  lineBuffer_6350 = _RAND_6357[7:0];
  _RAND_6358 = {1{`RANDOM}};
  lineBuffer_6351 = _RAND_6358[7:0];
  _RAND_6359 = {1{`RANDOM}};
  lineBuffer_6352 = _RAND_6359[7:0];
  _RAND_6360 = {1{`RANDOM}};
  lineBuffer_6353 = _RAND_6360[7:0];
  _RAND_6361 = {1{`RANDOM}};
  lineBuffer_6354 = _RAND_6361[7:0];
  _RAND_6362 = {1{`RANDOM}};
  lineBuffer_6355 = _RAND_6362[7:0];
  _RAND_6363 = {1{`RANDOM}};
  lineBuffer_6356 = _RAND_6363[7:0];
  _RAND_6364 = {1{`RANDOM}};
  lineBuffer_6357 = _RAND_6364[7:0];
  _RAND_6365 = {1{`RANDOM}};
  lineBuffer_6358 = _RAND_6365[7:0];
  _RAND_6366 = {1{`RANDOM}};
  lineBuffer_6359 = _RAND_6366[7:0];
  _RAND_6367 = {1{`RANDOM}};
  lineBuffer_6360 = _RAND_6367[7:0];
  _RAND_6368 = {1{`RANDOM}};
  lineBuffer_6361 = _RAND_6368[7:0];
  _RAND_6369 = {1{`RANDOM}};
  lineBuffer_6362 = _RAND_6369[7:0];
  _RAND_6370 = {1{`RANDOM}};
  lineBuffer_6363 = _RAND_6370[7:0];
  _RAND_6371 = {1{`RANDOM}};
  lineBuffer_6364 = _RAND_6371[7:0];
  _RAND_6372 = {1{`RANDOM}};
  lineBuffer_6365 = _RAND_6372[7:0];
  _RAND_6373 = {1{`RANDOM}};
  lineBuffer_6366 = _RAND_6373[7:0];
  _RAND_6374 = {1{`RANDOM}};
  lineBuffer_6367 = _RAND_6374[7:0];
  _RAND_6375 = {1{`RANDOM}};
  lineBuffer_6368 = _RAND_6375[7:0];
  _RAND_6376 = {1{`RANDOM}};
  lineBuffer_6369 = _RAND_6376[7:0];
  _RAND_6377 = {1{`RANDOM}};
  lineBuffer_6370 = _RAND_6377[7:0];
  _RAND_6378 = {1{`RANDOM}};
  lineBuffer_6371 = _RAND_6378[7:0];
  _RAND_6379 = {1{`RANDOM}};
  lineBuffer_6372 = _RAND_6379[7:0];
  _RAND_6380 = {1{`RANDOM}};
  lineBuffer_6373 = _RAND_6380[7:0];
  _RAND_6381 = {1{`RANDOM}};
  lineBuffer_6374 = _RAND_6381[7:0];
  _RAND_6382 = {1{`RANDOM}};
  lineBuffer_6375 = _RAND_6382[7:0];
  _RAND_6383 = {1{`RANDOM}};
  lineBuffer_6376 = _RAND_6383[7:0];
  _RAND_6384 = {1{`RANDOM}};
  lineBuffer_6377 = _RAND_6384[7:0];
  _RAND_6385 = {1{`RANDOM}};
  lineBuffer_6378 = _RAND_6385[7:0];
  _RAND_6386 = {1{`RANDOM}};
  lineBuffer_6379 = _RAND_6386[7:0];
  _RAND_6387 = {1{`RANDOM}};
  lineBuffer_6380 = _RAND_6387[7:0];
  _RAND_6388 = {1{`RANDOM}};
  lineBuffer_6381 = _RAND_6388[7:0];
  _RAND_6389 = {1{`RANDOM}};
  lineBuffer_6382 = _RAND_6389[7:0];
  _RAND_6390 = {1{`RANDOM}};
  lineBuffer_6383 = _RAND_6390[7:0];
  _RAND_6391 = {1{`RANDOM}};
  lineBuffer_6384 = _RAND_6391[7:0];
  _RAND_6392 = {1{`RANDOM}};
  lineBuffer_6385 = _RAND_6392[7:0];
  _RAND_6393 = {1{`RANDOM}};
  lineBuffer_6386 = _RAND_6393[7:0];
  _RAND_6394 = {1{`RANDOM}};
  lineBuffer_6387 = _RAND_6394[7:0];
  _RAND_6395 = {1{`RANDOM}};
  lineBuffer_6388 = _RAND_6395[7:0];
  _RAND_6396 = {1{`RANDOM}};
  lineBuffer_6389 = _RAND_6396[7:0];
  _RAND_6397 = {1{`RANDOM}};
  lineBuffer_6390 = _RAND_6397[7:0];
  _RAND_6398 = {1{`RANDOM}};
  lineBuffer_6391 = _RAND_6398[7:0];
  _RAND_6399 = {1{`RANDOM}};
  lineBuffer_6392 = _RAND_6399[7:0];
  _RAND_6400 = {1{`RANDOM}};
  lineBuffer_6393 = _RAND_6400[7:0];
  _RAND_6401 = {1{`RANDOM}};
  lineBuffer_6394 = _RAND_6401[7:0];
  _RAND_6402 = {1{`RANDOM}};
  lineBuffer_6395 = _RAND_6402[7:0];
  _RAND_6403 = {1{`RANDOM}};
  lineBuffer_6396 = _RAND_6403[7:0];
  _RAND_6404 = {1{`RANDOM}};
  lineBuffer_6397 = _RAND_6404[7:0];
  _RAND_6405 = {1{`RANDOM}};
  lineBuffer_6398 = _RAND_6405[7:0];
  _RAND_6406 = {1{`RANDOM}};
  lineBuffer_6399 = _RAND_6406[7:0];
  _RAND_6407 = {1{`RANDOM}};
  windowBuffer_0 = _RAND_6407[7:0];
  _RAND_6408 = {1{`RANDOM}};
  windowBuffer_1 = _RAND_6408[7:0];
  _RAND_6409 = {1{`RANDOM}};
  windowBuffer_2 = _RAND_6409[7:0];
  _RAND_6410 = {1{`RANDOM}};
  windowBuffer_3 = _RAND_6410[7:0];
  _RAND_6411 = {1{`RANDOM}};
  windowBuffer_4 = _RAND_6411[7:0];
  _RAND_6412 = {1{`RANDOM}};
  windowBuffer_5 = _RAND_6412[7:0];
  _RAND_6413 = {1{`RANDOM}};
  windowBuffer_6 = _RAND_6413[7:0];
  _RAND_6414 = {1{`RANDOM}};
  windowBuffer_7 = _RAND_6414[7:0];
  _RAND_6415 = {1{`RANDOM}};
  windowBuffer_8 = _RAND_6415[7:0];
  _RAND_6416 = {1{`RANDOM}};
  windowBuffer_9 = _RAND_6416[7:0];
  _RAND_6417 = {1{`RANDOM}};
  windowBuffer_10 = _RAND_6417[7:0];
  _RAND_6418 = {1{`RANDOM}};
  windowBuffer_11 = _RAND_6418[7:0];
  _RAND_6419 = {1{`RANDOM}};
  windowBuffer_12 = _RAND_6419[7:0];
  _RAND_6420 = {1{`RANDOM}};
  windowBuffer_13 = _RAND_6420[7:0];
  _RAND_6421 = {1{`RANDOM}};
  windowBuffer_14 = _RAND_6421[7:0];
  _RAND_6422 = {1{`RANDOM}};
  windowBuffer_15 = _RAND_6422[7:0];
  _RAND_6423 = {1{`RANDOM}};
  windowBuffer_16 = _RAND_6423[7:0];
  _RAND_6424 = {1{`RANDOM}};
  windowBuffer_17 = _RAND_6424[7:0];
  _RAND_6425 = {1{`RANDOM}};
  windowBuffer_18 = _RAND_6425[7:0];
  _RAND_6426 = {1{`RANDOM}};
  windowBuffer_19 = _RAND_6426[7:0];
  _RAND_6427 = {1{`RANDOM}};
  windowBuffer_20 = _RAND_6427[7:0];
  _RAND_6428 = {1{`RANDOM}};
  windowBuffer_21 = _RAND_6428[7:0];
  _RAND_6429 = {1{`RANDOM}};
  windowBuffer_22 = _RAND_6429[7:0];
  _RAND_6430 = {1{`RANDOM}};
  windowBuffer_23 = _RAND_6430[7:0];
  _RAND_6431 = {1{`RANDOM}};
  windowBuffer_24 = _RAND_6431[7:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      stateReg <= 2'h0;
    end else if (_T) begin
      if (io_enq_valid) begin
        stateReg <= 2'h1;
      end
    end else if (_T_1) begin
      if (_T_3) begin
        stateReg <= 2'h0;
      end else if (_T_4) begin
        stateReg <= 2'h1;
      end else if (_T_6) begin
        stateReg <= 2'h2;
      end
    end else if (_T_7) begin
      if (io_deq_ready) begin
        stateReg <= 2'h1;
      end
    end else if (_T_8) begin
      stateReg <= 2'h0;
    end
    if (_T) begin
      if (io_enq_valid) begin
        dataReg <= io_enq_bits;
      end
    end else if (_T_1) begin
      if (!(_T_3)) begin
        if (_T_4) begin
          dataReg <= io_enq_bits;
        end
      end
    end else if (_T_7) begin
      if (io_deq_ready) begin
        dataReg <= shadowReg;
      end
    end
    if (!(_T)) begin
      if (_T_1) begin
        if (!(_T_3)) begin
          if (!(_T_4)) begin
            if (_T_6) begin
              shadowReg <= io_enq_bits;
            end
          end
        end
      end
    end
    if (_T) begin
      userReg <= io_enq_user;
    end else if (_T_1) begin
      if (_T_3) begin
        userReg <= io_enq_user;
      end else if (_T_4) begin
        userReg <= io_enq_user;
      end
    end else if (_T_7) begin
      if (io_deq_ready) begin
        userReg <= shadowUserReg;
      end
    end
    if (!(_T)) begin
      if (_T_1) begin
        if (!(_T_3)) begin
          if (!(_T_4)) begin
            if (_T_6) begin
              shadowUserReg <= io_enq_user;
            end
          end
        end
      end
    end
    if (_T) begin
      if (io_enq_valid) begin
        lastReg <= io_enq_last;
      end
    end else if (_T_1) begin
      if (!(_T_3)) begin
        if (_T_4) begin
          lastReg <= io_enq_last;
        end
      end
    end else if (_T_7) begin
      if (io_deq_ready) begin
        lastReg <= shadowLastReg;
      end
    end
    if (!(_T)) begin
      if (_T_1) begin
        if (!(_T_3)) begin
          if (!(_T_4)) begin
            if (_T_6) begin
              shadowLastReg <= io_enq_last;
            end
          end
        end
      end
    end
    if (sel) begin
      lineBuffer_0 <= dataReg;
    end
    if (sel) begin
      lineBuffer_1 <= lineBuffer_0;
    end
    if (sel) begin
      lineBuffer_2 <= lineBuffer_1;
    end
    if (sel) begin
      lineBuffer_3 <= lineBuffer_2;
    end
    if (sel) begin
      lineBuffer_4 <= lineBuffer_3;
    end
    if (sel) begin
      lineBuffer_5 <= lineBuffer_4;
    end
    if (sel) begin
      lineBuffer_6 <= lineBuffer_5;
    end
    if (sel) begin
      lineBuffer_7 <= lineBuffer_6;
    end
    if (sel) begin
      lineBuffer_8 <= lineBuffer_7;
    end
    if (sel) begin
      lineBuffer_9 <= lineBuffer_8;
    end
    if (sel) begin
      lineBuffer_10 <= lineBuffer_9;
    end
    if (sel) begin
      lineBuffer_11 <= lineBuffer_10;
    end
    if (sel) begin
      lineBuffer_12 <= lineBuffer_11;
    end
    if (sel) begin
      lineBuffer_13 <= lineBuffer_12;
    end
    if (sel) begin
      lineBuffer_14 <= lineBuffer_13;
    end
    if (sel) begin
      lineBuffer_15 <= lineBuffer_14;
    end
    if (sel) begin
      lineBuffer_16 <= lineBuffer_15;
    end
    if (sel) begin
      lineBuffer_17 <= lineBuffer_16;
    end
    if (sel) begin
      lineBuffer_18 <= lineBuffer_17;
    end
    if (sel) begin
      lineBuffer_19 <= lineBuffer_18;
    end
    if (sel) begin
      lineBuffer_20 <= lineBuffer_19;
    end
    if (sel) begin
      lineBuffer_21 <= lineBuffer_20;
    end
    if (sel) begin
      lineBuffer_22 <= lineBuffer_21;
    end
    if (sel) begin
      lineBuffer_23 <= lineBuffer_22;
    end
    if (sel) begin
      lineBuffer_24 <= lineBuffer_23;
    end
    if (sel) begin
      lineBuffer_25 <= lineBuffer_24;
    end
    if (sel) begin
      lineBuffer_26 <= lineBuffer_25;
    end
    if (sel) begin
      lineBuffer_27 <= lineBuffer_26;
    end
    if (sel) begin
      lineBuffer_28 <= lineBuffer_27;
    end
    if (sel) begin
      lineBuffer_29 <= lineBuffer_28;
    end
    if (sel) begin
      lineBuffer_30 <= lineBuffer_29;
    end
    if (sel) begin
      lineBuffer_31 <= lineBuffer_30;
    end
    if (sel) begin
      lineBuffer_32 <= lineBuffer_31;
    end
    if (sel) begin
      lineBuffer_33 <= lineBuffer_32;
    end
    if (sel) begin
      lineBuffer_34 <= lineBuffer_33;
    end
    if (sel) begin
      lineBuffer_35 <= lineBuffer_34;
    end
    if (sel) begin
      lineBuffer_36 <= lineBuffer_35;
    end
    if (sel) begin
      lineBuffer_37 <= lineBuffer_36;
    end
    if (sel) begin
      lineBuffer_38 <= lineBuffer_37;
    end
    if (sel) begin
      lineBuffer_39 <= lineBuffer_38;
    end
    if (sel) begin
      lineBuffer_40 <= lineBuffer_39;
    end
    if (sel) begin
      lineBuffer_41 <= lineBuffer_40;
    end
    if (sel) begin
      lineBuffer_42 <= lineBuffer_41;
    end
    if (sel) begin
      lineBuffer_43 <= lineBuffer_42;
    end
    if (sel) begin
      lineBuffer_44 <= lineBuffer_43;
    end
    if (sel) begin
      lineBuffer_45 <= lineBuffer_44;
    end
    if (sel) begin
      lineBuffer_46 <= lineBuffer_45;
    end
    if (sel) begin
      lineBuffer_47 <= lineBuffer_46;
    end
    if (sel) begin
      lineBuffer_48 <= lineBuffer_47;
    end
    if (sel) begin
      lineBuffer_49 <= lineBuffer_48;
    end
    if (sel) begin
      lineBuffer_50 <= lineBuffer_49;
    end
    if (sel) begin
      lineBuffer_51 <= lineBuffer_50;
    end
    if (sel) begin
      lineBuffer_52 <= lineBuffer_51;
    end
    if (sel) begin
      lineBuffer_53 <= lineBuffer_52;
    end
    if (sel) begin
      lineBuffer_54 <= lineBuffer_53;
    end
    if (sel) begin
      lineBuffer_55 <= lineBuffer_54;
    end
    if (sel) begin
      lineBuffer_56 <= lineBuffer_55;
    end
    if (sel) begin
      lineBuffer_57 <= lineBuffer_56;
    end
    if (sel) begin
      lineBuffer_58 <= lineBuffer_57;
    end
    if (sel) begin
      lineBuffer_59 <= lineBuffer_58;
    end
    if (sel) begin
      lineBuffer_60 <= lineBuffer_59;
    end
    if (sel) begin
      lineBuffer_61 <= lineBuffer_60;
    end
    if (sel) begin
      lineBuffer_62 <= lineBuffer_61;
    end
    if (sel) begin
      lineBuffer_63 <= lineBuffer_62;
    end
    if (sel) begin
      lineBuffer_64 <= lineBuffer_63;
    end
    if (sel) begin
      lineBuffer_65 <= lineBuffer_64;
    end
    if (sel) begin
      lineBuffer_66 <= lineBuffer_65;
    end
    if (sel) begin
      lineBuffer_67 <= lineBuffer_66;
    end
    if (sel) begin
      lineBuffer_68 <= lineBuffer_67;
    end
    if (sel) begin
      lineBuffer_69 <= lineBuffer_68;
    end
    if (sel) begin
      lineBuffer_70 <= lineBuffer_69;
    end
    if (sel) begin
      lineBuffer_71 <= lineBuffer_70;
    end
    if (sel) begin
      lineBuffer_72 <= lineBuffer_71;
    end
    if (sel) begin
      lineBuffer_73 <= lineBuffer_72;
    end
    if (sel) begin
      lineBuffer_74 <= lineBuffer_73;
    end
    if (sel) begin
      lineBuffer_75 <= lineBuffer_74;
    end
    if (sel) begin
      lineBuffer_76 <= lineBuffer_75;
    end
    if (sel) begin
      lineBuffer_77 <= lineBuffer_76;
    end
    if (sel) begin
      lineBuffer_78 <= lineBuffer_77;
    end
    if (sel) begin
      lineBuffer_79 <= lineBuffer_78;
    end
    if (sel) begin
      lineBuffer_80 <= lineBuffer_79;
    end
    if (sel) begin
      lineBuffer_81 <= lineBuffer_80;
    end
    if (sel) begin
      lineBuffer_82 <= lineBuffer_81;
    end
    if (sel) begin
      lineBuffer_83 <= lineBuffer_82;
    end
    if (sel) begin
      lineBuffer_84 <= lineBuffer_83;
    end
    if (sel) begin
      lineBuffer_85 <= lineBuffer_84;
    end
    if (sel) begin
      lineBuffer_86 <= lineBuffer_85;
    end
    if (sel) begin
      lineBuffer_87 <= lineBuffer_86;
    end
    if (sel) begin
      lineBuffer_88 <= lineBuffer_87;
    end
    if (sel) begin
      lineBuffer_89 <= lineBuffer_88;
    end
    if (sel) begin
      lineBuffer_90 <= lineBuffer_89;
    end
    if (sel) begin
      lineBuffer_91 <= lineBuffer_90;
    end
    if (sel) begin
      lineBuffer_92 <= lineBuffer_91;
    end
    if (sel) begin
      lineBuffer_93 <= lineBuffer_92;
    end
    if (sel) begin
      lineBuffer_94 <= lineBuffer_93;
    end
    if (sel) begin
      lineBuffer_95 <= lineBuffer_94;
    end
    if (sel) begin
      lineBuffer_96 <= lineBuffer_95;
    end
    if (sel) begin
      lineBuffer_97 <= lineBuffer_96;
    end
    if (sel) begin
      lineBuffer_98 <= lineBuffer_97;
    end
    if (sel) begin
      lineBuffer_99 <= lineBuffer_98;
    end
    if (sel) begin
      lineBuffer_100 <= lineBuffer_99;
    end
    if (sel) begin
      lineBuffer_101 <= lineBuffer_100;
    end
    if (sel) begin
      lineBuffer_102 <= lineBuffer_101;
    end
    if (sel) begin
      lineBuffer_103 <= lineBuffer_102;
    end
    if (sel) begin
      lineBuffer_104 <= lineBuffer_103;
    end
    if (sel) begin
      lineBuffer_105 <= lineBuffer_104;
    end
    if (sel) begin
      lineBuffer_106 <= lineBuffer_105;
    end
    if (sel) begin
      lineBuffer_107 <= lineBuffer_106;
    end
    if (sel) begin
      lineBuffer_108 <= lineBuffer_107;
    end
    if (sel) begin
      lineBuffer_109 <= lineBuffer_108;
    end
    if (sel) begin
      lineBuffer_110 <= lineBuffer_109;
    end
    if (sel) begin
      lineBuffer_111 <= lineBuffer_110;
    end
    if (sel) begin
      lineBuffer_112 <= lineBuffer_111;
    end
    if (sel) begin
      lineBuffer_113 <= lineBuffer_112;
    end
    if (sel) begin
      lineBuffer_114 <= lineBuffer_113;
    end
    if (sel) begin
      lineBuffer_115 <= lineBuffer_114;
    end
    if (sel) begin
      lineBuffer_116 <= lineBuffer_115;
    end
    if (sel) begin
      lineBuffer_117 <= lineBuffer_116;
    end
    if (sel) begin
      lineBuffer_118 <= lineBuffer_117;
    end
    if (sel) begin
      lineBuffer_119 <= lineBuffer_118;
    end
    if (sel) begin
      lineBuffer_120 <= lineBuffer_119;
    end
    if (sel) begin
      lineBuffer_121 <= lineBuffer_120;
    end
    if (sel) begin
      lineBuffer_122 <= lineBuffer_121;
    end
    if (sel) begin
      lineBuffer_123 <= lineBuffer_122;
    end
    if (sel) begin
      lineBuffer_124 <= lineBuffer_123;
    end
    if (sel) begin
      lineBuffer_125 <= lineBuffer_124;
    end
    if (sel) begin
      lineBuffer_126 <= lineBuffer_125;
    end
    if (sel) begin
      lineBuffer_127 <= lineBuffer_126;
    end
    if (sel) begin
      lineBuffer_128 <= lineBuffer_127;
    end
    if (sel) begin
      lineBuffer_129 <= lineBuffer_128;
    end
    if (sel) begin
      lineBuffer_130 <= lineBuffer_129;
    end
    if (sel) begin
      lineBuffer_131 <= lineBuffer_130;
    end
    if (sel) begin
      lineBuffer_132 <= lineBuffer_131;
    end
    if (sel) begin
      lineBuffer_133 <= lineBuffer_132;
    end
    if (sel) begin
      lineBuffer_134 <= lineBuffer_133;
    end
    if (sel) begin
      lineBuffer_135 <= lineBuffer_134;
    end
    if (sel) begin
      lineBuffer_136 <= lineBuffer_135;
    end
    if (sel) begin
      lineBuffer_137 <= lineBuffer_136;
    end
    if (sel) begin
      lineBuffer_138 <= lineBuffer_137;
    end
    if (sel) begin
      lineBuffer_139 <= lineBuffer_138;
    end
    if (sel) begin
      lineBuffer_140 <= lineBuffer_139;
    end
    if (sel) begin
      lineBuffer_141 <= lineBuffer_140;
    end
    if (sel) begin
      lineBuffer_142 <= lineBuffer_141;
    end
    if (sel) begin
      lineBuffer_143 <= lineBuffer_142;
    end
    if (sel) begin
      lineBuffer_144 <= lineBuffer_143;
    end
    if (sel) begin
      lineBuffer_145 <= lineBuffer_144;
    end
    if (sel) begin
      lineBuffer_146 <= lineBuffer_145;
    end
    if (sel) begin
      lineBuffer_147 <= lineBuffer_146;
    end
    if (sel) begin
      lineBuffer_148 <= lineBuffer_147;
    end
    if (sel) begin
      lineBuffer_149 <= lineBuffer_148;
    end
    if (sel) begin
      lineBuffer_150 <= lineBuffer_149;
    end
    if (sel) begin
      lineBuffer_151 <= lineBuffer_150;
    end
    if (sel) begin
      lineBuffer_152 <= lineBuffer_151;
    end
    if (sel) begin
      lineBuffer_153 <= lineBuffer_152;
    end
    if (sel) begin
      lineBuffer_154 <= lineBuffer_153;
    end
    if (sel) begin
      lineBuffer_155 <= lineBuffer_154;
    end
    if (sel) begin
      lineBuffer_156 <= lineBuffer_155;
    end
    if (sel) begin
      lineBuffer_157 <= lineBuffer_156;
    end
    if (sel) begin
      lineBuffer_158 <= lineBuffer_157;
    end
    if (sel) begin
      lineBuffer_159 <= lineBuffer_158;
    end
    if (sel) begin
      lineBuffer_160 <= lineBuffer_159;
    end
    if (sel) begin
      lineBuffer_161 <= lineBuffer_160;
    end
    if (sel) begin
      lineBuffer_162 <= lineBuffer_161;
    end
    if (sel) begin
      lineBuffer_163 <= lineBuffer_162;
    end
    if (sel) begin
      lineBuffer_164 <= lineBuffer_163;
    end
    if (sel) begin
      lineBuffer_165 <= lineBuffer_164;
    end
    if (sel) begin
      lineBuffer_166 <= lineBuffer_165;
    end
    if (sel) begin
      lineBuffer_167 <= lineBuffer_166;
    end
    if (sel) begin
      lineBuffer_168 <= lineBuffer_167;
    end
    if (sel) begin
      lineBuffer_169 <= lineBuffer_168;
    end
    if (sel) begin
      lineBuffer_170 <= lineBuffer_169;
    end
    if (sel) begin
      lineBuffer_171 <= lineBuffer_170;
    end
    if (sel) begin
      lineBuffer_172 <= lineBuffer_171;
    end
    if (sel) begin
      lineBuffer_173 <= lineBuffer_172;
    end
    if (sel) begin
      lineBuffer_174 <= lineBuffer_173;
    end
    if (sel) begin
      lineBuffer_175 <= lineBuffer_174;
    end
    if (sel) begin
      lineBuffer_176 <= lineBuffer_175;
    end
    if (sel) begin
      lineBuffer_177 <= lineBuffer_176;
    end
    if (sel) begin
      lineBuffer_178 <= lineBuffer_177;
    end
    if (sel) begin
      lineBuffer_179 <= lineBuffer_178;
    end
    if (sel) begin
      lineBuffer_180 <= lineBuffer_179;
    end
    if (sel) begin
      lineBuffer_181 <= lineBuffer_180;
    end
    if (sel) begin
      lineBuffer_182 <= lineBuffer_181;
    end
    if (sel) begin
      lineBuffer_183 <= lineBuffer_182;
    end
    if (sel) begin
      lineBuffer_184 <= lineBuffer_183;
    end
    if (sel) begin
      lineBuffer_185 <= lineBuffer_184;
    end
    if (sel) begin
      lineBuffer_186 <= lineBuffer_185;
    end
    if (sel) begin
      lineBuffer_187 <= lineBuffer_186;
    end
    if (sel) begin
      lineBuffer_188 <= lineBuffer_187;
    end
    if (sel) begin
      lineBuffer_189 <= lineBuffer_188;
    end
    if (sel) begin
      lineBuffer_190 <= lineBuffer_189;
    end
    if (sel) begin
      lineBuffer_191 <= lineBuffer_190;
    end
    if (sel) begin
      lineBuffer_192 <= lineBuffer_191;
    end
    if (sel) begin
      lineBuffer_193 <= lineBuffer_192;
    end
    if (sel) begin
      lineBuffer_194 <= lineBuffer_193;
    end
    if (sel) begin
      lineBuffer_195 <= lineBuffer_194;
    end
    if (sel) begin
      lineBuffer_196 <= lineBuffer_195;
    end
    if (sel) begin
      lineBuffer_197 <= lineBuffer_196;
    end
    if (sel) begin
      lineBuffer_198 <= lineBuffer_197;
    end
    if (sel) begin
      lineBuffer_199 <= lineBuffer_198;
    end
    if (sel) begin
      lineBuffer_200 <= lineBuffer_199;
    end
    if (sel) begin
      lineBuffer_201 <= lineBuffer_200;
    end
    if (sel) begin
      lineBuffer_202 <= lineBuffer_201;
    end
    if (sel) begin
      lineBuffer_203 <= lineBuffer_202;
    end
    if (sel) begin
      lineBuffer_204 <= lineBuffer_203;
    end
    if (sel) begin
      lineBuffer_205 <= lineBuffer_204;
    end
    if (sel) begin
      lineBuffer_206 <= lineBuffer_205;
    end
    if (sel) begin
      lineBuffer_207 <= lineBuffer_206;
    end
    if (sel) begin
      lineBuffer_208 <= lineBuffer_207;
    end
    if (sel) begin
      lineBuffer_209 <= lineBuffer_208;
    end
    if (sel) begin
      lineBuffer_210 <= lineBuffer_209;
    end
    if (sel) begin
      lineBuffer_211 <= lineBuffer_210;
    end
    if (sel) begin
      lineBuffer_212 <= lineBuffer_211;
    end
    if (sel) begin
      lineBuffer_213 <= lineBuffer_212;
    end
    if (sel) begin
      lineBuffer_214 <= lineBuffer_213;
    end
    if (sel) begin
      lineBuffer_215 <= lineBuffer_214;
    end
    if (sel) begin
      lineBuffer_216 <= lineBuffer_215;
    end
    if (sel) begin
      lineBuffer_217 <= lineBuffer_216;
    end
    if (sel) begin
      lineBuffer_218 <= lineBuffer_217;
    end
    if (sel) begin
      lineBuffer_219 <= lineBuffer_218;
    end
    if (sel) begin
      lineBuffer_220 <= lineBuffer_219;
    end
    if (sel) begin
      lineBuffer_221 <= lineBuffer_220;
    end
    if (sel) begin
      lineBuffer_222 <= lineBuffer_221;
    end
    if (sel) begin
      lineBuffer_223 <= lineBuffer_222;
    end
    if (sel) begin
      lineBuffer_224 <= lineBuffer_223;
    end
    if (sel) begin
      lineBuffer_225 <= lineBuffer_224;
    end
    if (sel) begin
      lineBuffer_226 <= lineBuffer_225;
    end
    if (sel) begin
      lineBuffer_227 <= lineBuffer_226;
    end
    if (sel) begin
      lineBuffer_228 <= lineBuffer_227;
    end
    if (sel) begin
      lineBuffer_229 <= lineBuffer_228;
    end
    if (sel) begin
      lineBuffer_230 <= lineBuffer_229;
    end
    if (sel) begin
      lineBuffer_231 <= lineBuffer_230;
    end
    if (sel) begin
      lineBuffer_232 <= lineBuffer_231;
    end
    if (sel) begin
      lineBuffer_233 <= lineBuffer_232;
    end
    if (sel) begin
      lineBuffer_234 <= lineBuffer_233;
    end
    if (sel) begin
      lineBuffer_235 <= lineBuffer_234;
    end
    if (sel) begin
      lineBuffer_236 <= lineBuffer_235;
    end
    if (sel) begin
      lineBuffer_237 <= lineBuffer_236;
    end
    if (sel) begin
      lineBuffer_238 <= lineBuffer_237;
    end
    if (sel) begin
      lineBuffer_239 <= lineBuffer_238;
    end
    if (sel) begin
      lineBuffer_240 <= lineBuffer_239;
    end
    if (sel) begin
      lineBuffer_241 <= lineBuffer_240;
    end
    if (sel) begin
      lineBuffer_242 <= lineBuffer_241;
    end
    if (sel) begin
      lineBuffer_243 <= lineBuffer_242;
    end
    if (sel) begin
      lineBuffer_244 <= lineBuffer_243;
    end
    if (sel) begin
      lineBuffer_245 <= lineBuffer_244;
    end
    if (sel) begin
      lineBuffer_246 <= lineBuffer_245;
    end
    if (sel) begin
      lineBuffer_247 <= lineBuffer_246;
    end
    if (sel) begin
      lineBuffer_248 <= lineBuffer_247;
    end
    if (sel) begin
      lineBuffer_249 <= lineBuffer_248;
    end
    if (sel) begin
      lineBuffer_250 <= lineBuffer_249;
    end
    if (sel) begin
      lineBuffer_251 <= lineBuffer_250;
    end
    if (sel) begin
      lineBuffer_252 <= lineBuffer_251;
    end
    if (sel) begin
      lineBuffer_253 <= lineBuffer_252;
    end
    if (sel) begin
      lineBuffer_254 <= lineBuffer_253;
    end
    if (sel) begin
      lineBuffer_255 <= lineBuffer_254;
    end
    if (sel) begin
      lineBuffer_256 <= lineBuffer_255;
    end
    if (sel) begin
      lineBuffer_257 <= lineBuffer_256;
    end
    if (sel) begin
      lineBuffer_258 <= lineBuffer_257;
    end
    if (sel) begin
      lineBuffer_259 <= lineBuffer_258;
    end
    if (sel) begin
      lineBuffer_260 <= lineBuffer_259;
    end
    if (sel) begin
      lineBuffer_261 <= lineBuffer_260;
    end
    if (sel) begin
      lineBuffer_262 <= lineBuffer_261;
    end
    if (sel) begin
      lineBuffer_263 <= lineBuffer_262;
    end
    if (sel) begin
      lineBuffer_264 <= lineBuffer_263;
    end
    if (sel) begin
      lineBuffer_265 <= lineBuffer_264;
    end
    if (sel) begin
      lineBuffer_266 <= lineBuffer_265;
    end
    if (sel) begin
      lineBuffer_267 <= lineBuffer_266;
    end
    if (sel) begin
      lineBuffer_268 <= lineBuffer_267;
    end
    if (sel) begin
      lineBuffer_269 <= lineBuffer_268;
    end
    if (sel) begin
      lineBuffer_270 <= lineBuffer_269;
    end
    if (sel) begin
      lineBuffer_271 <= lineBuffer_270;
    end
    if (sel) begin
      lineBuffer_272 <= lineBuffer_271;
    end
    if (sel) begin
      lineBuffer_273 <= lineBuffer_272;
    end
    if (sel) begin
      lineBuffer_274 <= lineBuffer_273;
    end
    if (sel) begin
      lineBuffer_275 <= lineBuffer_274;
    end
    if (sel) begin
      lineBuffer_276 <= lineBuffer_275;
    end
    if (sel) begin
      lineBuffer_277 <= lineBuffer_276;
    end
    if (sel) begin
      lineBuffer_278 <= lineBuffer_277;
    end
    if (sel) begin
      lineBuffer_279 <= lineBuffer_278;
    end
    if (sel) begin
      lineBuffer_280 <= lineBuffer_279;
    end
    if (sel) begin
      lineBuffer_281 <= lineBuffer_280;
    end
    if (sel) begin
      lineBuffer_282 <= lineBuffer_281;
    end
    if (sel) begin
      lineBuffer_283 <= lineBuffer_282;
    end
    if (sel) begin
      lineBuffer_284 <= lineBuffer_283;
    end
    if (sel) begin
      lineBuffer_285 <= lineBuffer_284;
    end
    if (sel) begin
      lineBuffer_286 <= lineBuffer_285;
    end
    if (sel) begin
      lineBuffer_287 <= lineBuffer_286;
    end
    if (sel) begin
      lineBuffer_288 <= lineBuffer_287;
    end
    if (sel) begin
      lineBuffer_289 <= lineBuffer_288;
    end
    if (sel) begin
      lineBuffer_290 <= lineBuffer_289;
    end
    if (sel) begin
      lineBuffer_291 <= lineBuffer_290;
    end
    if (sel) begin
      lineBuffer_292 <= lineBuffer_291;
    end
    if (sel) begin
      lineBuffer_293 <= lineBuffer_292;
    end
    if (sel) begin
      lineBuffer_294 <= lineBuffer_293;
    end
    if (sel) begin
      lineBuffer_295 <= lineBuffer_294;
    end
    if (sel) begin
      lineBuffer_296 <= lineBuffer_295;
    end
    if (sel) begin
      lineBuffer_297 <= lineBuffer_296;
    end
    if (sel) begin
      lineBuffer_298 <= lineBuffer_297;
    end
    if (sel) begin
      lineBuffer_299 <= lineBuffer_298;
    end
    if (sel) begin
      lineBuffer_300 <= lineBuffer_299;
    end
    if (sel) begin
      lineBuffer_301 <= lineBuffer_300;
    end
    if (sel) begin
      lineBuffer_302 <= lineBuffer_301;
    end
    if (sel) begin
      lineBuffer_303 <= lineBuffer_302;
    end
    if (sel) begin
      lineBuffer_304 <= lineBuffer_303;
    end
    if (sel) begin
      lineBuffer_305 <= lineBuffer_304;
    end
    if (sel) begin
      lineBuffer_306 <= lineBuffer_305;
    end
    if (sel) begin
      lineBuffer_307 <= lineBuffer_306;
    end
    if (sel) begin
      lineBuffer_308 <= lineBuffer_307;
    end
    if (sel) begin
      lineBuffer_309 <= lineBuffer_308;
    end
    if (sel) begin
      lineBuffer_310 <= lineBuffer_309;
    end
    if (sel) begin
      lineBuffer_311 <= lineBuffer_310;
    end
    if (sel) begin
      lineBuffer_312 <= lineBuffer_311;
    end
    if (sel) begin
      lineBuffer_313 <= lineBuffer_312;
    end
    if (sel) begin
      lineBuffer_314 <= lineBuffer_313;
    end
    if (sel) begin
      lineBuffer_315 <= lineBuffer_314;
    end
    if (sel) begin
      lineBuffer_316 <= lineBuffer_315;
    end
    if (sel) begin
      lineBuffer_317 <= lineBuffer_316;
    end
    if (sel) begin
      lineBuffer_318 <= lineBuffer_317;
    end
    if (sel) begin
      lineBuffer_319 <= lineBuffer_318;
    end
    if (sel) begin
      lineBuffer_320 <= lineBuffer_319;
    end
    if (sel) begin
      lineBuffer_321 <= lineBuffer_320;
    end
    if (sel) begin
      lineBuffer_322 <= lineBuffer_321;
    end
    if (sel) begin
      lineBuffer_323 <= lineBuffer_322;
    end
    if (sel) begin
      lineBuffer_324 <= lineBuffer_323;
    end
    if (sel) begin
      lineBuffer_325 <= lineBuffer_324;
    end
    if (sel) begin
      lineBuffer_326 <= lineBuffer_325;
    end
    if (sel) begin
      lineBuffer_327 <= lineBuffer_326;
    end
    if (sel) begin
      lineBuffer_328 <= lineBuffer_327;
    end
    if (sel) begin
      lineBuffer_329 <= lineBuffer_328;
    end
    if (sel) begin
      lineBuffer_330 <= lineBuffer_329;
    end
    if (sel) begin
      lineBuffer_331 <= lineBuffer_330;
    end
    if (sel) begin
      lineBuffer_332 <= lineBuffer_331;
    end
    if (sel) begin
      lineBuffer_333 <= lineBuffer_332;
    end
    if (sel) begin
      lineBuffer_334 <= lineBuffer_333;
    end
    if (sel) begin
      lineBuffer_335 <= lineBuffer_334;
    end
    if (sel) begin
      lineBuffer_336 <= lineBuffer_335;
    end
    if (sel) begin
      lineBuffer_337 <= lineBuffer_336;
    end
    if (sel) begin
      lineBuffer_338 <= lineBuffer_337;
    end
    if (sel) begin
      lineBuffer_339 <= lineBuffer_338;
    end
    if (sel) begin
      lineBuffer_340 <= lineBuffer_339;
    end
    if (sel) begin
      lineBuffer_341 <= lineBuffer_340;
    end
    if (sel) begin
      lineBuffer_342 <= lineBuffer_341;
    end
    if (sel) begin
      lineBuffer_343 <= lineBuffer_342;
    end
    if (sel) begin
      lineBuffer_344 <= lineBuffer_343;
    end
    if (sel) begin
      lineBuffer_345 <= lineBuffer_344;
    end
    if (sel) begin
      lineBuffer_346 <= lineBuffer_345;
    end
    if (sel) begin
      lineBuffer_347 <= lineBuffer_346;
    end
    if (sel) begin
      lineBuffer_348 <= lineBuffer_347;
    end
    if (sel) begin
      lineBuffer_349 <= lineBuffer_348;
    end
    if (sel) begin
      lineBuffer_350 <= lineBuffer_349;
    end
    if (sel) begin
      lineBuffer_351 <= lineBuffer_350;
    end
    if (sel) begin
      lineBuffer_352 <= lineBuffer_351;
    end
    if (sel) begin
      lineBuffer_353 <= lineBuffer_352;
    end
    if (sel) begin
      lineBuffer_354 <= lineBuffer_353;
    end
    if (sel) begin
      lineBuffer_355 <= lineBuffer_354;
    end
    if (sel) begin
      lineBuffer_356 <= lineBuffer_355;
    end
    if (sel) begin
      lineBuffer_357 <= lineBuffer_356;
    end
    if (sel) begin
      lineBuffer_358 <= lineBuffer_357;
    end
    if (sel) begin
      lineBuffer_359 <= lineBuffer_358;
    end
    if (sel) begin
      lineBuffer_360 <= lineBuffer_359;
    end
    if (sel) begin
      lineBuffer_361 <= lineBuffer_360;
    end
    if (sel) begin
      lineBuffer_362 <= lineBuffer_361;
    end
    if (sel) begin
      lineBuffer_363 <= lineBuffer_362;
    end
    if (sel) begin
      lineBuffer_364 <= lineBuffer_363;
    end
    if (sel) begin
      lineBuffer_365 <= lineBuffer_364;
    end
    if (sel) begin
      lineBuffer_366 <= lineBuffer_365;
    end
    if (sel) begin
      lineBuffer_367 <= lineBuffer_366;
    end
    if (sel) begin
      lineBuffer_368 <= lineBuffer_367;
    end
    if (sel) begin
      lineBuffer_369 <= lineBuffer_368;
    end
    if (sel) begin
      lineBuffer_370 <= lineBuffer_369;
    end
    if (sel) begin
      lineBuffer_371 <= lineBuffer_370;
    end
    if (sel) begin
      lineBuffer_372 <= lineBuffer_371;
    end
    if (sel) begin
      lineBuffer_373 <= lineBuffer_372;
    end
    if (sel) begin
      lineBuffer_374 <= lineBuffer_373;
    end
    if (sel) begin
      lineBuffer_375 <= lineBuffer_374;
    end
    if (sel) begin
      lineBuffer_376 <= lineBuffer_375;
    end
    if (sel) begin
      lineBuffer_377 <= lineBuffer_376;
    end
    if (sel) begin
      lineBuffer_378 <= lineBuffer_377;
    end
    if (sel) begin
      lineBuffer_379 <= lineBuffer_378;
    end
    if (sel) begin
      lineBuffer_380 <= lineBuffer_379;
    end
    if (sel) begin
      lineBuffer_381 <= lineBuffer_380;
    end
    if (sel) begin
      lineBuffer_382 <= lineBuffer_381;
    end
    if (sel) begin
      lineBuffer_383 <= lineBuffer_382;
    end
    if (sel) begin
      lineBuffer_384 <= lineBuffer_383;
    end
    if (sel) begin
      lineBuffer_385 <= lineBuffer_384;
    end
    if (sel) begin
      lineBuffer_386 <= lineBuffer_385;
    end
    if (sel) begin
      lineBuffer_387 <= lineBuffer_386;
    end
    if (sel) begin
      lineBuffer_388 <= lineBuffer_387;
    end
    if (sel) begin
      lineBuffer_389 <= lineBuffer_388;
    end
    if (sel) begin
      lineBuffer_390 <= lineBuffer_389;
    end
    if (sel) begin
      lineBuffer_391 <= lineBuffer_390;
    end
    if (sel) begin
      lineBuffer_392 <= lineBuffer_391;
    end
    if (sel) begin
      lineBuffer_393 <= lineBuffer_392;
    end
    if (sel) begin
      lineBuffer_394 <= lineBuffer_393;
    end
    if (sel) begin
      lineBuffer_395 <= lineBuffer_394;
    end
    if (sel) begin
      lineBuffer_396 <= lineBuffer_395;
    end
    if (sel) begin
      lineBuffer_397 <= lineBuffer_396;
    end
    if (sel) begin
      lineBuffer_398 <= lineBuffer_397;
    end
    if (sel) begin
      lineBuffer_399 <= lineBuffer_398;
    end
    if (sel) begin
      lineBuffer_400 <= lineBuffer_399;
    end
    if (sel) begin
      lineBuffer_401 <= lineBuffer_400;
    end
    if (sel) begin
      lineBuffer_402 <= lineBuffer_401;
    end
    if (sel) begin
      lineBuffer_403 <= lineBuffer_402;
    end
    if (sel) begin
      lineBuffer_404 <= lineBuffer_403;
    end
    if (sel) begin
      lineBuffer_405 <= lineBuffer_404;
    end
    if (sel) begin
      lineBuffer_406 <= lineBuffer_405;
    end
    if (sel) begin
      lineBuffer_407 <= lineBuffer_406;
    end
    if (sel) begin
      lineBuffer_408 <= lineBuffer_407;
    end
    if (sel) begin
      lineBuffer_409 <= lineBuffer_408;
    end
    if (sel) begin
      lineBuffer_410 <= lineBuffer_409;
    end
    if (sel) begin
      lineBuffer_411 <= lineBuffer_410;
    end
    if (sel) begin
      lineBuffer_412 <= lineBuffer_411;
    end
    if (sel) begin
      lineBuffer_413 <= lineBuffer_412;
    end
    if (sel) begin
      lineBuffer_414 <= lineBuffer_413;
    end
    if (sel) begin
      lineBuffer_415 <= lineBuffer_414;
    end
    if (sel) begin
      lineBuffer_416 <= lineBuffer_415;
    end
    if (sel) begin
      lineBuffer_417 <= lineBuffer_416;
    end
    if (sel) begin
      lineBuffer_418 <= lineBuffer_417;
    end
    if (sel) begin
      lineBuffer_419 <= lineBuffer_418;
    end
    if (sel) begin
      lineBuffer_420 <= lineBuffer_419;
    end
    if (sel) begin
      lineBuffer_421 <= lineBuffer_420;
    end
    if (sel) begin
      lineBuffer_422 <= lineBuffer_421;
    end
    if (sel) begin
      lineBuffer_423 <= lineBuffer_422;
    end
    if (sel) begin
      lineBuffer_424 <= lineBuffer_423;
    end
    if (sel) begin
      lineBuffer_425 <= lineBuffer_424;
    end
    if (sel) begin
      lineBuffer_426 <= lineBuffer_425;
    end
    if (sel) begin
      lineBuffer_427 <= lineBuffer_426;
    end
    if (sel) begin
      lineBuffer_428 <= lineBuffer_427;
    end
    if (sel) begin
      lineBuffer_429 <= lineBuffer_428;
    end
    if (sel) begin
      lineBuffer_430 <= lineBuffer_429;
    end
    if (sel) begin
      lineBuffer_431 <= lineBuffer_430;
    end
    if (sel) begin
      lineBuffer_432 <= lineBuffer_431;
    end
    if (sel) begin
      lineBuffer_433 <= lineBuffer_432;
    end
    if (sel) begin
      lineBuffer_434 <= lineBuffer_433;
    end
    if (sel) begin
      lineBuffer_435 <= lineBuffer_434;
    end
    if (sel) begin
      lineBuffer_436 <= lineBuffer_435;
    end
    if (sel) begin
      lineBuffer_437 <= lineBuffer_436;
    end
    if (sel) begin
      lineBuffer_438 <= lineBuffer_437;
    end
    if (sel) begin
      lineBuffer_439 <= lineBuffer_438;
    end
    if (sel) begin
      lineBuffer_440 <= lineBuffer_439;
    end
    if (sel) begin
      lineBuffer_441 <= lineBuffer_440;
    end
    if (sel) begin
      lineBuffer_442 <= lineBuffer_441;
    end
    if (sel) begin
      lineBuffer_443 <= lineBuffer_442;
    end
    if (sel) begin
      lineBuffer_444 <= lineBuffer_443;
    end
    if (sel) begin
      lineBuffer_445 <= lineBuffer_444;
    end
    if (sel) begin
      lineBuffer_446 <= lineBuffer_445;
    end
    if (sel) begin
      lineBuffer_447 <= lineBuffer_446;
    end
    if (sel) begin
      lineBuffer_448 <= lineBuffer_447;
    end
    if (sel) begin
      lineBuffer_449 <= lineBuffer_448;
    end
    if (sel) begin
      lineBuffer_450 <= lineBuffer_449;
    end
    if (sel) begin
      lineBuffer_451 <= lineBuffer_450;
    end
    if (sel) begin
      lineBuffer_452 <= lineBuffer_451;
    end
    if (sel) begin
      lineBuffer_453 <= lineBuffer_452;
    end
    if (sel) begin
      lineBuffer_454 <= lineBuffer_453;
    end
    if (sel) begin
      lineBuffer_455 <= lineBuffer_454;
    end
    if (sel) begin
      lineBuffer_456 <= lineBuffer_455;
    end
    if (sel) begin
      lineBuffer_457 <= lineBuffer_456;
    end
    if (sel) begin
      lineBuffer_458 <= lineBuffer_457;
    end
    if (sel) begin
      lineBuffer_459 <= lineBuffer_458;
    end
    if (sel) begin
      lineBuffer_460 <= lineBuffer_459;
    end
    if (sel) begin
      lineBuffer_461 <= lineBuffer_460;
    end
    if (sel) begin
      lineBuffer_462 <= lineBuffer_461;
    end
    if (sel) begin
      lineBuffer_463 <= lineBuffer_462;
    end
    if (sel) begin
      lineBuffer_464 <= lineBuffer_463;
    end
    if (sel) begin
      lineBuffer_465 <= lineBuffer_464;
    end
    if (sel) begin
      lineBuffer_466 <= lineBuffer_465;
    end
    if (sel) begin
      lineBuffer_467 <= lineBuffer_466;
    end
    if (sel) begin
      lineBuffer_468 <= lineBuffer_467;
    end
    if (sel) begin
      lineBuffer_469 <= lineBuffer_468;
    end
    if (sel) begin
      lineBuffer_470 <= lineBuffer_469;
    end
    if (sel) begin
      lineBuffer_471 <= lineBuffer_470;
    end
    if (sel) begin
      lineBuffer_472 <= lineBuffer_471;
    end
    if (sel) begin
      lineBuffer_473 <= lineBuffer_472;
    end
    if (sel) begin
      lineBuffer_474 <= lineBuffer_473;
    end
    if (sel) begin
      lineBuffer_475 <= lineBuffer_474;
    end
    if (sel) begin
      lineBuffer_476 <= lineBuffer_475;
    end
    if (sel) begin
      lineBuffer_477 <= lineBuffer_476;
    end
    if (sel) begin
      lineBuffer_478 <= lineBuffer_477;
    end
    if (sel) begin
      lineBuffer_479 <= lineBuffer_478;
    end
    if (sel) begin
      lineBuffer_480 <= lineBuffer_479;
    end
    if (sel) begin
      lineBuffer_481 <= lineBuffer_480;
    end
    if (sel) begin
      lineBuffer_482 <= lineBuffer_481;
    end
    if (sel) begin
      lineBuffer_483 <= lineBuffer_482;
    end
    if (sel) begin
      lineBuffer_484 <= lineBuffer_483;
    end
    if (sel) begin
      lineBuffer_485 <= lineBuffer_484;
    end
    if (sel) begin
      lineBuffer_486 <= lineBuffer_485;
    end
    if (sel) begin
      lineBuffer_487 <= lineBuffer_486;
    end
    if (sel) begin
      lineBuffer_488 <= lineBuffer_487;
    end
    if (sel) begin
      lineBuffer_489 <= lineBuffer_488;
    end
    if (sel) begin
      lineBuffer_490 <= lineBuffer_489;
    end
    if (sel) begin
      lineBuffer_491 <= lineBuffer_490;
    end
    if (sel) begin
      lineBuffer_492 <= lineBuffer_491;
    end
    if (sel) begin
      lineBuffer_493 <= lineBuffer_492;
    end
    if (sel) begin
      lineBuffer_494 <= lineBuffer_493;
    end
    if (sel) begin
      lineBuffer_495 <= lineBuffer_494;
    end
    if (sel) begin
      lineBuffer_496 <= lineBuffer_495;
    end
    if (sel) begin
      lineBuffer_497 <= lineBuffer_496;
    end
    if (sel) begin
      lineBuffer_498 <= lineBuffer_497;
    end
    if (sel) begin
      lineBuffer_499 <= lineBuffer_498;
    end
    if (sel) begin
      lineBuffer_500 <= lineBuffer_499;
    end
    if (sel) begin
      lineBuffer_501 <= lineBuffer_500;
    end
    if (sel) begin
      lineBuffer_502 <= lineBuffer_501;
    end
    if (sel) begin
      lineBuffer_503 <= lineBuffer_502;
    end
    if (sel) begin
      lineBuffer_504 <= lineBuffer_503;
    end
    if (sel) begin
      lineBuffer_505 <= lineBuffer_504;
    end
    if (sel) begin
      lineBuffer_506 <= lineBuffer_505;
    end
    if (sel) begin
      lineBuffer_507 <= lineBuffer_506;
    end
    if (sel) begin
      lineBuffer_508 <= lineBuffer_507;
    end
    if (sel) begin
      lineBuffer_509 <= lineBuffer_508;
    end
    if (sel) begin
      lineBuffer_510 <= lineBuffer_509;
    end
    if (sel) begin
      lineBuffer_511 <= lineBuffer_510;
    end
    if (sel) begin
      lineBuffer_512 <= lineBuffer_511;
    end
    if (sel) begin
      lineBuffer_513 <= lineBuffer_512;
    end
    if (sel) begin
      lineBuffer_514 <= lineBuffer_513;
    end
    if (sel) begin
      lineBuffer_515 <= lineBuffer_514;
    end
    if (sel) begin
      lineBuffer_516 <= lineBuffer_515;
    end
    if (sel) begin
      lineBuffer_517 <= lineBuffer_516;
    end
    if (sel) begin
      lineBuffer_518 <= lineBuffer_517;
    end
    if (sel) begin
      lineBuffer_519 <= lineBuffer_518;
    end
    if (sel) begin
      lineBuffer_520 <= lineBuffer_519;
    end
    if (sel) begin
      lineBuffer_521 <= lineBuffer_520;
    end
    if (sel) begin
      lineBuffer_522 <= lineBuffer_521;
    end
    if (sel) begin
      lineBuffer_523 <= lineBuffer_522;
    end
    if (sel) begin
      lineBuffer_524 <= lineBuffer_523;
    end
    if (sel) begin
      lineBuffer_525 <= lineBuffer_524;
    end
    if (sel) begin
      lineBuffer_526 <= lineBuffer_525;
    end
    if (sel) begin
      lineBuffer_527 <= lineBuffer_526;
    end
    if (sel) begin
      lineBuffer_528 <= lineBuffer_527;
    end
    if (sel) begin
      lineBuffer_529 <= lineBuffer_528;
    end
    if (sel) begin
      lineBuffer_530 <= lineBuffer_529;
    end
    if (sel) begin
      lineBuffer_531 <= lineBuffer_530;
    end
    if (sel) begin
      lineBuffer_532 <= lineBuffer_531;
    end
    if (sel) begin
      lineBuffer_533 <= lineBuffer_532;
    end
    if (sel) begin
      lineBuffer_534 <= lineBuffer_533;
    end
    if (sel) begin
      lineBuffer_535 <= lineBuffer_534;
    end
    if (sel) begin
      lineBuffer_536 <= lineBuffer_535;
    end
    if (sel) begin
      lineBuffer_537 <= lineBuffer_536;
    end
    if (sel) begin
      lineBuffer_538 <= lineBuffer_537;
    end
    if (sel) begin
      lineBuffer_539 <= lineBuffer_538;
    end
    if (sel) begin
      lineBuffer_540 <= lineBuffer_539;
    end
    if (sel) begin
      lineBuffer_541 <= lineBuffer_540;
    end
    if (sel) begin
      lineBuffer_542 <= lineBuffer_541;
    end
    if (sel) begin
      lineBuffer_543 <= lineBuffer_542;
    end
    if (sel) begin
      lineBuffer_544 <= lineBuffer_543;
    end
    if (sel) begin
      lineBuffer_545 <= lineBuffer_544;
    end
    if (sel) begin
      lineBuffer_546 <= lineBuffer_545;
    end
    if (sel) begin
      lineBuffer_547 <= lineBuffer_546;
    end
    if (sel) begin
      lineBuffer_548 <= lineBuffer_547;
    end
    if (sel) begin
      lineBuffer_549 <= lineBuffer_548;
    end
    if (sel) begin
      lineBuffer_550 <= lineBuffer_549;
    end
    if (sel) begin
      lineBuffer_551 <= lineBuffer_550;
    end
    if (sel) begin
      lineBuffer_552 <= lineBuffer_551;
    end
    if (sel) begin
      lineBuffer_553 <= lineBuffer_552;
    end
    if (sel) begin
      lineBuffer_554 <= lineBuffer_553;
    end
    if (sel) begin
      lineBuffer_555 <= lineBuffer_554;
    end
    if (sel) begin
      lineBuffer_556 <= lineBuffer_555;
    end
    if (sel) begin
      lineBuffer_557 <= lineBuffer_556;
    end
    if (sel) begin
      lineBuffer_558 <= lineBuffer_557;
    end
    if (sel) begin
      lineBuffer_559 <= lineBuffer_558;
    end
    if (sel) begin
      lineBuffer_560 <= lineBuffer_559;
    end
    if (sel) begin
      lineBuffer_561 <= lineBuffer_560;
    end
    if (sel) begin
      lineBuffer_562 <= lineBuffer_561;
    end
    if (sel) begin
      lineBuffer_563 <= lineBuffer_562;
    end
    if (sel) begin
      lineBuffer_564 <= lineBuffer_563;
    end
    if (sel) begin
      lineBuffer_565 <= lineBuffer_564;
    end
    if (sel) begin
      lineBuffer_566 <= lineBuffer_565;
    end
    if (sel) begin
      lineBuffer_567 <= lineBuffer_566;
    end
    if (sel) begin
      lineBuffer_568 <= lineBuffer_567;
    end
    if (sel) begin
      lineBuffer_569 <= lineBuffer_568;
    end
    if (sel) begin
      lineBuffer_570 <= lineBuffer_569;
    end
    if (sel) begin
      lineBuffer_571 <= lineBuffer_570;
    end
    if (sel) begin
      lineBuffer_572 <= lineBuffer_571;
    end
    if (sel) begin
      lineBuffer_573 <= lineBuffer_572;
    end
    if (sel) begin
      lineBuffer_574 <= lineBuffer_573;
    end
    if (sel) begin
      lineBuffer_575 <= lineBuffer_574;
    end
    if (sel) begin
      lineBuffer_576 <= lineBuffer_575;
    end
    if (sel) begin
      lineBuffer_577 <= lineBuffer_576;
    end
    if (sel) begin
      lineBuffer_578 <= lineBuffer_577;
    end
    if (sel) begin
      lineBuffer_579 <= lineBuffer_578;
    end
    if (sel) begin
      lineBuffer_580 <= lineBuffer_579;
    end
    if (sel) begin
      lineBuffer_581 <= lineBuffer_580;
    end
    if (sel) begin
      lineBuffer_582 <= lineBuffer_581;
    end
    if (sel) begin
      lineBuffer_583 <= lineBuffer_582;
    end
    if (sel) begin
      lineBuffer_584 <= lineBuffer_583;
    end
    if (sel) begin
      lineBuffer_585 <= lineBuffer_584;
    end
    if (sel) begin
      lineBuffer_586 <= lineBuffer_585;
    end
    if (sel) begin
      lineBuffer_587 <= lineBuffer_586;
    end
    if (sel) begin
      lineBuffer_588 <= lineBuffer_587;
    end
    if (sel) begin
      lineBuffer_589 <= lineBuffer_588;
    end
    if (sel) begin
      lineBuffer_590 <= lineBuffer_589;
    end
    if (sel) begin
      lineBuffer_591 <= lineBuffer_590;
    end
    if (sel) begin
      lineBuffer_592 <= lineBuffer_591;
    end
    if (sel) begin
      lineBuffer_593 <= lineBuffer_592;
    end
    if (sel) begin
      lineBuffer_594 <= lineBuffer_593;
    end
    if (sel) begin
      lineBuffer_595 <= lineBuffer_594;
    end
    if (sel) begin
      lineBuffer_596 <= lineBuffer_595;
    end
    if (sel) begin
      lineBuffer_597 <= lineBuffer_596;
    end
    if (sel) begin
      lineBuffer_598 <= lineBuffer_597;
    end
    if (sel) begin
      lineBuffer_599 <= lineBuffer_598;
    end
    if (sel) begin
      lineBuffer_600 <= lineBuffer_599;
    end
    if (sel) begin
      lineBuffer_601 <= lineBuffer_600;
    end
    if (sel) begin
      lineBuffer_602 <= lineBuffer_601;
    end
    if (sel) begin
      lineBuffer_603 <= lineBuffer_602;
    end
    if (sel) begin
      lineBuffer_604 <= lineBuffer_603;
    end
    if (sel) begin
      lineBuffer_605 <= lineBuffer_604;
    end
    if (sel) begin
      lineBuffer_606 <= lineBuffer_605;
    end
    if (sel) begin
      lineBuffer_607 <= lineBuffer_606;
    end
    if (sel) begin
      lineBuffer_608 <= lineBuffer_607;
    end
    if (sel) begin
      lineBuffer_609 <= lineBuffer_608;
    end
    if (sel) begin
      lineBuffer_610 <= lineBuffer_609;
    end
    if (sel) begin
      lineBuffer_611 <= lineBuffer_610;
    end
    if (sel) begin
      lineBuffer_612 <= lineBuffer_611;
    end
    if (sel) begin
      lineBuffer_613 <= lineBuffer_612;
    end
    if (sel) begin
      lineBuffer_614 <= lineBuffer_613;
    end
    if (sel) begin
      lineBuffer_615 <= lineBuffer_614;
    end
    if (sel) begin
      lineBuffer_616 <= lineBuffer_615;
    end
    if (sel) begin
      lineBuffer_617 <= lineBuffer_616;
    end
    if (sel) begin
      lineBuffer_618 <= lineBuffer_617;
    end
    if (sel) begin
      lineBuffer_619 <= lineBuffer_618;
    end
    if (sel) begin
      lineBuffer_620 <= lineBuffer_619;
    end
    if (sel) begin
      lineBuffer_621 <= lineBuffer_620;
    end
    if (sel) begin
      lineBuffer_622 <= lineBuffer_621;
    end
    if (sel) begin
      lineBuffer_623 <= lineBuffer_622;
    end
    if (sel) begin
      lineBuffer_624 <= lineBuffer_623;
    end
    if (sel) begin
      lineBuffer_625 <= lineBuffer_624;
    end
    if (sel) begin
      lineBuffer_626 <= lineBuffer_625;
    end
    if (sel) begin
      lineBuffer_627 <= lineBuffer_626;
    end
    if (sel) begin
      lineBuffer_628 <= lineBuffer_627;
    end
    if (sel) begin
      lineBuffer_629 <= lineBuffer_628;
    end
    if (sel) begin
      lineBuffer_630 <= lineBuffer_629;
    end
    if (sel) begin
      lineBuffer_631 <= lineBuffer_630;
    end
    if (sel) begin
      lineBuffer_632 <= lineBuffer_631;
    end
    if (sel) begin
      lineBuffer_633 <= lineBuffer_632;
    end
    if (sel) begin
      lineBuffer_634 <= lineBuffer_633;
    end
    if (sel) begin
      lineBuffer_635 <= lineBuffer_634;
    end
    if (sel) begin
      lineBuffer_636 <= lineBuffer_635;
    end
    if (sel) begin
      lineBuffer_637 <= lineBuffer_636;
    end
    if (sel) begin
      lineBuffer_638 <= lineBuffer_637;
    end
    if (sel) begin
      lineBuffer_639 <= lineBuffer_638;
    end
    if (sel) begin
      lineBuffer_640 <= lineBuffer_639;
    end
    if (sel) begin
      lineBuffer_641 <= lineBuffer_640;
    end
    if (sel) begin
      lineBuffer_642 <= lineBuffer_641;
    end
    if (sel) begin
      lineBuffer_643 <= lineBuffer_642;
    end
    if (sel) begin
      lineBuffer_644 <= lineBuffer_643;
    end
    if (sel) begin
      lineBuffer_645 <= lineBuffer_644;
    end
    if (sel) begin
      lineBuffer_646 <= lineBuffer_645;
    end
    if (sel) begin
      lineBuffer_647 <= lineBuffer_646;
    end
    if (sel) begin
      lineBuffer_648 <= lineBuffer_647;
    end
    if (sel) begin
      lineBuffer_649 <= lineBuffer_648;
    end
    if (sel) begin
      lineBuffer_650 <= lineBuffer_649;
    end
    if (sel) begin
      lineBuffer_651 <= lineBuffer_650;
    end
    if (sel) begin
      lineBuffer_652 <= lineBuffer_651;
    end
    if (sel) begin
      lineBuffer_653 <= lineBuffer_652;
    end
    if (sel) begin
      lineBuffer_654 <= lineBuffer_653;
    end
    if (sel) begin
      lineBuffer_655 <= lineBuffer_654;
    end
    if (sel) begin
      lineBuffer_656 <= lineBuffer_655;
    end
    if (sel) begin
      lineBuffer_657 <= lineBuffer_656;
    end
    if (sel) begin
      lineBuffer_658 <= lineBuffer_657;
    end
    if (sel) begin
      lineBuffer_659 <= lineBuffer_658;
    end
    if (sel) begin
      lineBuffer_660 <= lineBuffer_659;
    end
    if (sel) begin
      lineBuffer_661 <= lineBuffer_660;
    end
    if (sel) begin
      lineBuffer_662 <= lineBuffer_661;
    end
    if (sel) begin
      lineBuffer_663 <= lineBuffer_662;
    end
    if (sel) begin
      lineBuffer_664 <= lineBuffer_663;
    end
    if (sel) begin
      lineBuffer_665 <= lineBuffer_664;
    end
    if (sel) begin
      lineBuffer_666 <= lineBuffer_665;
    end
    if (sel) begin
      lineBuffer_667 <= lineBuffer_666;
    end
    if (sel) begin
      lineBuffer_668 <= lineBuffer_667;
    end
    if (sel) begin
      lineBuffer_669 <= lineBuffer_668;
    end
    if (sel) begin
      lineBuffer_670 <= lineBuffer_669;
    end
    if (sel) begin
      lineBuffer_671 <= lineBuffer_670;
    end
    if (sel) begin
      lineBuffer_672 <= lineBuffer_671;
    end
    if (sel) begin
      lineBuffer_673 <= lineBuffer_672;
    end
    if (sel) begin
      lineBuffer_674 <= lineBuffer_673;
    end
    if (sel) begin
      lineBuffer_675 <= lineBuffer_674;
    end
    if (sel) begin
      lineBuffer_676 <= lineBuffer_675;
    end
    if (sel) begin
      lineBuffer_677 <= lineBuffer_676;
    end
    if (sel) begin
      lineBuffer_678 <= lineBuffer_677;
    end
    if (sel) begin
      lineBuffer_679 <= lineBuffer_678;
    end
    if (sel) begin
      lineBuffer_680 <= lineBuffer_679;
    end
    if (sel) begin
      lineBuffer_681 <= lineBuffer_680;
    end
    if (sel) begin
      lineBuffer_682 <= lineBuffer_681;
    end
    if (sel) begin
      lineBuffer_683 <= lineBuffer_682;
    end
    if (sel) begin
      lineBuffer_684 <= lineBuffer_683;
    end
    if (sel) begin
      lineBuffer_685 <= lineBuffer_684;
    end
    if (sel) begin
      lineBuffer_686 <= lineBuffer_685;
    end
    if (sel) begin
      lineBuffer_687 <= lineBuffer_686;
    end
    if (sel) begin
      lineBuffer_688 <= lineBuffer_687;
    end
    if (sel) begin
      lineBuffer_689 <= lineBuffer_688;
    end
    if (sel) begin
      lineBuffer_690 <= lineBuffer_689;
    end
    if (sel) begin
      lineBuffer_691 <= lineBuffer_690;
    end
    if (sel) begin
      lineBuffer_692 <= lineBuffer_691;
    end
    if (sel) begin
      lineBuffer_693 <= lineBuffer_692;
    end
    if (sel) begin
      lineBuffer_694 <= lineBuffer_693;
    end
    if (sel) begin
      lineBuffer_695 <= lineBuffer_694;
    end
    if (sel) begin
      lineBuffer_696 <= lineBuffer_695;
    end
    if (sel) begin
      lineBuffer_697 <= lineBuffer_696;
    end
    if (sel) begin
      lineBuffer_698 <= lineBuffer_697;
    end
    if (sel) begin
      lineBuffer_699 <= lineBuffer_698;
    end
    if (sel) begin
      lineBuffer_700 <= lineBuffer_699;
    end
    if (sel) begin
      lineBuffer_701 <= lineBuffer_700;
    end
    if (sel) begin
      lineBuffer_702 <= lineBuffer_701;
    end
    if (sel) begin
      lineBuffer_703 <= lineBuffer_702;
    end
    if (sel) begin
      lineBuffer_704 <= lineBuffer_703;
    end
    if (sel) begin
      lineBuffer_705 <= lineBuffer_704;
    end
    if (sel) begin
      lineBuffer_706 <= lineBuffer_705;
    end
    if (sel) begin
      lineBuffer_707 <= lineBuffer_706;
    end
    if (sel) begin
      lineBuffer_708 <= lineBuffer_707;
    end
    if (sel) begin
      lineBuffer_709 <= lineBuffer_708;
    end
    if (sel) begin
      lineBuffer_710 <= lineBuffer_709;
    end
    if (sel) begin
      lineBuffer_711 <= lineBuffer_710;
    end
    if (sel) begin
      lineBuffer_712 <= lineBuffer_711;
    end
    if (sel) begin
      lineBuffer_713 <= lineBuffer_712;
    end
    if (sel) begin
      lineBuffer_714 <= lineBuffer_713;
    end
    if (sel) begin
      lineBuffer_715 <= lineBuffer_714;
    end
    if (sel) begin
      lineBuffer_716 <= lineBuffer_715;
    end
    if (sel) begin
      lineBuffer_717 <= lineBuffer_716;
    end
    if (sel) begin
      lineBuffer_718 <= lineBuffer_717;
    end
    if (sel) begin
      lineBuffer_719 <= lineBuffer_718;
    end
    if (sel) begin
      lineBuffer_720 <= lineBuffer_719;
    end
    if (sel) begin
      lineBuffer_721 <= lineBuffer_720;
    end
    if (sel) begin
      lineBuffer_722 <= lineBuffer_721;
    end
    if (sel) begin
      lineBuffer_723 <= lineBuffer_722;
    end
    if (sel) begin
      lineBuffer_724 <= lineBuffer_723;
    end
    if (sel) begin
      lineBuffer_725 <= lineBuffer_724;
    end
    if (sel) begin
      lineBuffer_726 <= lineBuffer_725;
    end
    if (sel) begin
      lineBuffer_727 <= lineBuffer_726;
    end
    if (sel) begin
      lineBuffer_728 <= lineBuffer_727;
    end
    if (sel) begin
      lineBuffer_729 <= lineBuffer_728;
    end
    if (sel) begin
      lineBuffer_730 <= lineBuffer_729;
    end
    if (sel) begin
      lineBuffer_731 <= lineBuffer_730;
    end
    if (sel) begin
      lineBuffer_732 <= lineBuffer_731;
    end
    if (sel) begin
      lineBuffer_733 <= lineBuffer_732;
    end
    if (sel) begin
      lineBuffer_734 <= lineBuffer_733;
    end
    if (sel) begin
      lineBuffer_735 <= lineBuffer_734;
    end
    if (sel) begin
      lineBuffer_736 <= lineBuffer_735;
    end
    if (sel) begin
      lineBuffer_737 <= lineBuffer_736;
    end
    if (sel) begin
      lineBuffer_738 <= lineBuffer_737;
    end
    if (sel) begin
      lineBuffer_739 <= lineBuffer_738;
    end
    if (sel) begin
      lineBuffer_740 <= lineBuffer_739;
    end
    if (sel) begin
      lineBuffer_741 <= lineBuffer_740;
    end
    if (sel) begin
      lineBuffer_742 <= lineBuffer_741;
    end
    if (sel) begin
      lineBuffer_743 <= lineBuffer_742;
    end
    if (sel) begin
      lineBuffer_744 <= lineBuffer_743;
    end
    if (sel) begin
      lineBuffer_745 <= lineBuffer_744;
    end
    if (sel) begin
      lineBuffer_746 <= lineBuffer_745;
    end
    if (sel) begin
      lineBuffer_747 <= lineBuffer_746;
    end
    if (sel) begin
      lineBuffer_748 <= lineBuffer_747;
    end
    if (sel) begin
      lineBuffer_749 <= lineBuffer_748;
    end
    if (sel) begin
      lineBuffer_750 <= lineBuffer_749;
    end
    if (sel) begin
      lineBuffer_751 <= lineBuffer_750;
    end
    if (sel) begin
      lineBuffer_752 <= lineBuffer_751;
    end
    if (sel) begin
      lineBuffer_753 <= lineBuffer_752;
    end
    if (sel) begin
      lineBuffer_754 <= lineBuffer_753;
    end
    if (sel) begin
      lineBuffer_755 <= lineBuffer_754;
    end
    if (sel) begin
      lineBuffer_756 <= lineBuffer_755;
    end
    if (sel) begin
      lineBuffer_757 <= lineBuffer_756;
    end
    if (sel) begin
      lineBuffer_758 <= lineBuffer_757;
    end
    if (sel) begin
      lineBuffer_759 <= lineBuffer_758;
    end
    if (sel) begin
      lineBuffer_760 <= lineBuffer_759;
    end
    if (sel) begin
      lineBuffer_761 <= lineBuffer_760;
    end
    if (sel) begin
      lineBuffer_762 <= lineBuffer_761;
    end
    if (sel) begin
      lineBuffer_763 <= lineBuffer_762;
    end
    if (sel) begin
      lineBuffer_764 <= lineBuffer_763;
    end
    if (sel) begin
      lineBuffer_765 <= lineBuffer_764;
    end
    if (sel) begin
      lineBuffer_766 <= lineBuffer_765;
    end
    if (sel) begin
      lineBuffer_767 <= lineBuffer_766;
    end
    if (sel) begin
      lineBuffer_768 <= lineBuffer_767;
    end
    if (sel) begin
      lineBuffer_769 <= lineBuffer_768;
    end
    if (sel) begin
      lineBuffer_770 <= lineBuffer_769;
    end
    if (sel) begin
      lineBuffer_771 <= lineBuffer_770;
    end
    if (sel) begin
      lineBuffer_772 <= lineBuffer_771;
    end
    if (sel) begin
      lineBuffer_773 <= lineBuffer_772;
    end
    if (sel) begin
      lineBuffer_774 <= lineBuffer_773;
    end
    if (sel) begin
      lineBuffer_775 <= lineBuffer_774;
    end
    if (sel) begin
      lineBuffer_776 <= lineBuffer_775;
    end
    if (sel) begin
      lineBuffer_777 <= lineBuffer_776;
    end
    if (sel) begin
      lineBuffer_778 <= lineBuffer_777;
    end
    if (sel) begin
      lineBuffer_779 <= lineBuffer_778;
    end
    if (sel) begin
      lineBuffer_780 <= lineBuffer_779;
    end
    if (sel) begin
      lineBuffer_781 <= lineBuffer_780;
    end
    if (sel) begin
      lineBuffer_782 <= lineBuffer_781;
    end
    if (sel) begin
      lineBuffer_783 <= lineBuffer_782;
    end
    if (sel) begin
      lineBuffer_784 <= lineBuffer_783;
    end
    if (sel) begin
      lineBuffer_785 <= lineBuffer_784;
    end
    if (sel) begin
      lineBuffer_786 <= lineBuffer_785;
    end
    if (sel) begin
      lineBuffer_787 <= lineBuffer_786;
    end
    if (sel) begin
      lineBuffer_788 <= lineBuffer_787;
    end
    if (sel) begin
      lineBuffer_789 <= lineBuffer_788;
    end
    if (sel) begin
      lineBuffer_790 <= lineBuffer_789;
    end
    if (sel) begin
      lineBuffer_791 <= lineBuffer_790;
    end
    if (sel) begin
      lineBuffer_792 <= lineBuffer_791;
    end
    if (sel) begin
      lineBuffer_793 <= lineBuffer_792;
    end
    if (sel) begin
      lineBuffer_794 <= lineBuffer_793;
    end
    if (sel) begin
      lineBuffer_795 <= lineBuffer_794;
    end
    if (sel) begin
      lineBuffer_796 <= lineBuffer_795;
    end
    if (sel) begin
      lineBuffer_797 <= lineBuffer_796;
    end
    if (sel) begin
      lineBuffer_798 <= lineBuffer_797;
    end
    if (sel) begin
      lineBuffer_799 <= lineBuffer_798;
    end
    if (sel) begin
      lineBuffer_800 <= lineBuffer_799;
    end
    if (sel) begin
      lineBuffer_801 <= lineBuffer_800;
    end
    if (sel) begin
      lineBuffer_802 <= lineBuffer_801;
    end
    if (sel) begin
      lineBuffer_803 <= lineBuffer_802;
    end
    if (sel) begin
      lineBuffer_804 <= lineBuffer_803;
    end
    if (sel) begin
      lineBuffer_805 <= lineBuffer_804;
    end
    if (sel) begin
      lineBuffer_806 <= lineBuffer_805;
    end
    if (sel) begin
      lineBuffer_807 <= lineBuffer_806;
    end
    if (sel) begin
      lineBuffer_808 <= lineBuffer_807;
    end
    if (sel) begin
      lineBuffer_809 <= lineBuffer_808;
    end
    if (sel) begin
      lineBuffer_810 <= lineBuffer_809;
    end
    if (sel) begin
      lineBuffer_811 <= lineBuffer_810;
    end
    if (sel) begin
      lineBuffer_812 <= lineBuffer_811;
    end
    if (sel) begin
      lineBuffer_813 <= lineBuffer_812;
    end
    if (sel) begin
      lineBuffer_814 <= lineBuffer_813;
    end
    if (sel) begin
      lineBuffer_815 <= lineBuffer_814;
    end
    if (sel) begin
      lineBuffer_816 <= lineBuffer_815;
    end
    if (sel) begin
      lineBuffer_817 <= lineBuffer_816;
    end
    if (sel) begin
      lineBuffer_818 <= lineBuffer_817;
    end
    if (sel) begin
      lineBuffer_819 <= lineBuffer_818;
    end
    if (sel) begin
      lineBuffer_820 <= lineBuffer_819;
    end
    if (sel) begin
      lineBuffer_821 <= lineBuffer_820;
    end
    if (sel) begin
      lineBuffer_822 <= lineBuffer_821;
    end
    if (sel) begin
      lineBuffer_823 <= lineBuffer_822;
    end
    if (sel) begin
      lineBuffer_824 <= lineBuffer_823;
    end
    if (sel) begin
      lineBuffer_825 <= lineBuffer_824;
    end
    if (sel) begin
      lineBuffer_826 <= lineBuffer_825;
    end
    if (sel) begin
      lineBuffer_827 <= lineBuffer_826;
    end
    if (sel) begin
      lineBuffer_828 <= lineBuffer_827;
    end
    if (sel) begin
      lineBuffer_829 <= lineBuffer_828;
    end
    if (sel) begin
      lineBuffer_830 <= lineBuffer_829;
    end
    if (sel) begin
      lineBuffer_831 <= lineBuffer_830;
    end
    if (sel) begin
      lineBuffer_832 <= lineBuffer_831;
    end
    if (sel) begin
      lineBuffer_833 <= lineBuffer_832;
    end
    if (sel) begin
      lineBuffer_834 <= lineBuffer_833;
    end
    if (sel) begin
      lineBuffer_835 <= lineBuffer_834;
    end
    if (sel) begin
      lineBuffer_836 <= lineBuffer_835;
    end
    if (sel) begin
      lineBuffer_837 <= lineBuffer_836;
    end
    if (sel) begin
      lineBuffer_838 <= lineBuffer_837;
    end
    if (sel) begin
      lineBuffer_839 <= lineBuffer_838;
    end
    if (sel) begin
      lineBuffer_840 <= lineBuffer_839;
    end
    if (sel) begin
      lineBuffer_841 <= lineBuffer_840;
    end
    if (sel) begin
      lineBuffer_842 <= lineBuffer_841;
    end
    if (sel) begin
      lineBuffer_843 <= lineBuffer_842;
    end
    if (sel) begin
      lineBuffer_844 <= lineBuffer_843;
    end
    if (sel) begin
      lineBuffer_845 <= lineBuffer_844;
    end
    if (sel) begin
      lineBuffer_846 <= lineBuffer_845;
    end
    if (sel) begin
      lineBuffer_847 <= lineBuffer_846;
    end
    if (sel) begin
      lineBuffer_848 <= lineBuffer_847;
    end
    if (sel) begin
      lineBuffer_849 <= lineBuffer_848;
    end
    if (sel) begin
      lineBuffer_850 <= lineBuffer_849;
    end
    if (sel) begin
      lineBuffer_851 <= lineBuffer_850;
    end
    if (sel) begin
      lineBuffer_852 <= lineBuffer_851;
    end
    if (sel) begin
      lineBuffer_853 <= lineBuffer_852;
    end
    if (sel) begin
      lineBuffer_854 <= lineBuffer_853;
    end
    if (sel) begin
      lineBuffer_855 <= lineBuffer_854;
    end
    if (sel) begin
      lineBuffer_856 <= lineBuffer_855;
    end
    if (sel) begin
      lineBuffer_857 <= lineBuffer_856;
    end
    if (sel) begin
      lineBuffer_858 <= lineBuffer_857;
    end
    if (sel) begin
      lineBuffer_859 <= lineBuffer_858;
    end
    if (sel) begin
      lineBuffer_860 <= lineBuffer_859;
    end
    if (sel) begin
      lineBuffer_861 <= lineBuffer_860;
    end
    if (sel) begin
      lineBuffer_862 <= lineBuffer_861;
    end
    if (sel) begin
      lineBuffer_863 <= lineBuffer_862;
    end
    if (sel) begin
      lineBuffer_864 <= lineBuffer_863;
    end
    if (sel) begin
      lineBuffer_865 <= lineBuffer_864;
    end
    if (sel) begin
      lineBuffer_866 <= lineBuffer_865;
    end
    if (sel) begin
      lineBuffer_867 <= lineBuffer_866;
    end
    if (sel) begin
      lineBuffer_868 <= lineBuffer_867;
    end
    if (sel) begin
      lineBuffer_869 <= lineBuffer_868;
    end
    if (sel) begin
      lineBuffer_870 <= lineBuffer_869;
    end
    if (sel) begin
      lineBuffer_871 <= lineBuffer_870;
    end
    if (sel) begin
      lineBuffer_872 <= lineBuffer_871;
    end
    if (sel) begin
      lineBuffer_873 <= lineBuffer_872;
    end
    if (sel) begin
      lineBuffer_874 <= lineBuffer_873;
    end
    if (sel) begin
      lineBuffer_875 <= lineBuffer_874;
    end
    if (sel) begin
      lineBuffer_876 <= lineBuffer_875;
    end
    if (sel) begin
      lineBuffer_877 <= lineBuffer_876;
    end
    if (sel) begin
      lineBuffer_878 <= lineBuffer_877;
    end
    if (sel) begin
      lineBuffer_879 <= lineBuffer_878;
    end
    if (sel) begin
      lineBuffer_880 <= lineBuffer_879;
    end
    if (sel) begin
      lineBuffer_881 <= lineBuffer_880;
    end
    if (sel) begin
      lineBuffer_882 <= lineBuffer_881;
    end
    if (sel) begin
      lineBuffer_883 <= lineBuffer_882;
    end
    if (sel) begin
      lineBuffer_884 <= lineBuffer_883;
    end
    if (sel) begin
      lineBuffer_885 <= lineBuffer_884;
    end
    if (sel) begin
      lineBuffer_886 <= lineBuffer_885;
    end
    if (sel) begin
      lineBuffer_887 <= lineBuffer_886;
    end
    if (sel) begin
      lineBuffer_888 <= lineBuffer_887;
    end
    if (sel) begin
      lineBuffer_889 <= lineBuffer_888;
    end
    if (sel) begin
      lineBuffer_890 <= lineBuffer_889;
    end
    if (sel) begin
      lineBuffer_891 <= lineBuffer_890;
    end
    if (sel) begin
      lineBuffer_892 <= lineBuffer_891;
    end
    if (sel) begin
      lineBuffer_893 <= lineBuffer_892;
    end
    if (sel) begin
      lineBuffer_894 <= lineBuffer_893;
    end
    if (sel) begin
      lineBuffer_895 <= lineBuffer_894;
    end
    if (sel) begin
      lineBuffer_896 <= lineBuffer_895;
    end
    if (sel) begin
      lineBuffer_897 <= lineBuffer_896;
    end
    if (sel) begin
      lineBuffer_898 <= lineBuffer_897;
    end
    if (sel) begin
      lineBuffer_899 <= lineBuffer_898;
    end
    if (sel) begin
      lineBuffer_900 <= lineBuffer_899;
    end
    if (sel) begin
      lineBuffer_901 <= lineBuffer_900;
    end
    if (sel) begin
      lineBuffer_902 <= lineBuffer_901;
    end
    if (sel) begin
      lineBuffer_903 <= lineBuffer_902;
    end
    if (sel) begin
      lineBuffer_904 <= lineBuffer_903;
    end
    if (sel) begin
      lineBuffer_905 <= lineBuffer_904;
    end
    if (sel) begin
      lineBuffer_906 <= lineBuffer_905;
    end
    if (sel) begin
      lineBuffer_907 <= lineBuffer_906;
    end
    if (sel) begin
      lineBuffer_908 <= lineBuffer_907;
    end
    if (sel) begin
      lineBuffer_909 <= lineBuffer_908;
    end
    if (sel) begin
      lineBuffer_910 <= lineBuffer_909;
    end
    if (sel) begin
      lineBuffer_911 <= lineBuffer_910;
    end
    if (sel) begin
      lineBuffer_912 <= lineBuffer_911;
    end
    if (sel) begin
      lineBuffer_913 <= lineBuffer_912;
    end
    if (sel) begin
      lineBuffer_914 <= lineBuffer_913;
    end
    if (sel) begin
      lineBuffer_915 <= lineBuffer_914;
    end
    if (sel) begin
      lineBuffer_916 <= lineBuffer_915;
    end
    if (sel) begin
      lineBuffer_917 <= lineBuffer_916;
    end
    if (sel) begin
      lineBuffer_918 <= lineBuffer_917;
    end
    if (sel) begin
      lineBuffer_919 <= lineBuffer_918;
    end
    if (sel) begin
      lineBuffer_920 <= lineBuffer_919;
    end
    if (sel) begin
      lineBuffer_921 <= lineBuffer_920;
    end
    if (sel) begin
      lineBuffer_922 <= lineBuffer_921;
    end
    if (sel) begin
      lineBuffer_923 <= lineBuffer_922;
    end
    if (sel) begin
      lineBuffer_924 <= lineBuffer_923;
    end
    if (sel) begin
      lineBuffer_925 <= lineBuffer_924;
    end
    if (sel) begin
      lineBuffer_926 <= lineBuffer_925;
    end
    if (sel) begin
      lineBuffer_927 <= lineBuffer_926;
    end
    if (sel) begin
      lineBuffer_928 <= lineBuffer_927;
    end
    if (sel) begin
      lineBuffer_929 <= lineBuffer_928;
    end
    if (sel) begin
      lineBuffer_930 <= lineBuffer_929;
    end
    if (sel) begin
      lineBuffer_931 <= lineBuffer_930;
    end
    if (sel) begin
      lineBuffer_932 <= lineBuffer_931;
    end
    if (sel) begin
      lineBuffer_933 <= lineBuffer_932;
    end
    if (sel) begin
      lineBuffer_934 <= lineBuffer_933;
    end
    if (sel) begin
      lineBuffer_935 <= lineBuffer_934;
    end
    if (sel) begin
      lineBuffer_936 <= lineBuffer_935;
    end
    if (sel) begin
      lineBuffer_937 <= lineBuffer_936;
    end
    if (sel) begin
      lineBuffer_938 <= lineBuffer_937;
    end
    if (sel) begin
      lineBuffer_939 <= lineBuffer_938;
    end
    if (sel) begin
      lineBuffer_940 <= lineBuffer_939;
    end
    if (sel) begin
      lineBuffer_941 <= lineBuffer_940;
    end
    if (sel) begin
      lineBuffer_942 <= lineBuffer_941;
    end
    if (sel) begin
      lineBuffer_943 <= lineBuffer_942;
    end
    if (sel) begin
      lineBuffer_944 <= lineBuffer_943;
    end
    if (sel) begin
      lineBuffer_945 <= lineBuffer_944;
    end
    if (sel) begin
      lineBuffer_946 <= lineBuffer_945;
    end
    if (sel) begin
      lineBuffer_947 <= lineBuffer_946;
    end
    if (sel) begin
      lineBuffer_948 <= lineBuffer_947;
    end
    if (sel) begin
      lineBuffer_949 <= lineBuffer_948;
    end
    if (sel) begin
      lineBuffer_950 <= lineBuffer_949;
    end
    if (sel) begin
      lineBuffer_951 <= lineBuffer_950;
    end
    if (sel) begin
      lineBuffer_952 <= lineBuffer_951;
    end
    if (sel) begin
      lineBuffer_953 <= lineBuffer_952;
    end
    if (sel) begin
      lineBuffer_954 <= lineBuffer_953;
    end
    if (sel) begin
      lineBuffer_955 <= lineBuffer_954;
    end
    if (sel) begin
      lineBuffer_956 <= lineBuffer_955;
    end
    if (sel) begin
      lineBuffer_957 <= lineBuffer_956;
    end
    if (sel) begin
      lineBuffer_958 <= lineBuffer_957;
    end
    if (sel) begin
      lineBuffer_959 <= lineBuffer_958;
    end
    if (sel) begin
      lineBuffer_960 <= lineBuffer_959;
    end
    if (sel) begin
      lineBuffer_961 <= lineBuffer_960;
    end
    if (sel) begin
      lineBuffer_962 <= lineBuffer_961;
    end
    if (sel) begin
      lineBuffer_963 <= lineBuffer_962;
    end
    if (sel) begin
      lineBuffer_964 <= lineBuffer_963;
    end
    if (sel) begin
      lineBuffer_965 <= lineBuffer_964;
    end
    if (sel) begin
      lineBuffer_966 <= lineBuffer_965;
    end
    if (sel) begin
      lineBuffer_967 <= lineBuffer_966;
    end
    if (sel) begin
      lineBuffer_968 <= lineBuffer_967;
    end
    if (sel) begin
      lineBuffer_969 <= lineBuffer_968;
    end
    if (sel) begin
      lineBuffer_970 <= lineBuffer_969;
    end
    if (sel) begin
      lineBuffer_971 <= lineBuffer_970;
    end
    if (sel) begin
      lineBuffer_972 <= lineBuffer_971;
    end
    if (sel) begin
      lineBuffer_973 <= lineBuffer_972;
    end
    if (sel) begin
      lineBuffer_974 <= lineBuffer_973;
    end
    if (sel) begin
      lineBuffer_975 <= lineBuffer_974;
    end
    if (sel) begin
      lineBuffer_976 <= lineBuffer_975;
    end
    if (sel) begin
      lineBuffer_977 <= lineBuffer_976;
    end
    if (sel) begin
      lineBuffer_978 <= lineBuffer_977;
    end
    if (sel) begin
      lineBuffer_979 <= lineBuffer_978;
    end
    if (sel) begin
      lineBuffer_980 <= lineBuffer_979;
    end
    if (sel) begin
      lineBuffer_981 <= lineBuffer_980;
    end
    if (sel) begin
      lineBuffer_982 <= lineBuffer_981;
    end
    if (sel) begin
      lineBuffer_983 <= lineBuffer_982;
    end
    if (sel) begin
      lineBuffer_984 <= lineBuffer_983;
    end
    if (sel) begin
      lineBuffer_985 <= lineBuffer_984;
    end
    if (sel) begin
      lineBuffer_986 <= lineBuffer_985;
    end
    if (sel) begin
      lineBuffer_987 <= lineBuffer_986;
    end
    if (sel) begin
      lineBuffer_988 <= lineBuffer_987;
    end
    if (sel) begin
      lineBuffer_989 <= lineBuffer_988;
    end
    if (sel) begin
      lineBuffer_990 <= lineBuffer_989;
    end
    if (sel) begin
      lineBuffer_991 <= lineBuffer_990;
    end
    if (sel) begin
      lineBuffer_992 <= lineBuffer_991;
    end
    if (sel) begin
      lineBuffer_993 <= lineBuffer_992;
    end
    if (sel) begin
      lineBuffer_994 <= lineBuffer_993;
    end
    if (sel) begin
      lineBuffer_995 <= lineBuffer_994;
    end
    if (sel) begin
      lineBuffer_996 <= lineBuffer_995;
    end
    if (sel) begin
      lineBuffer_997 <= lineBuffer_996;
    end
    if (sel) begin
      lineBuffer_998 <= lineBuffer_997;
    end
    if (sel) begin
      lineBuffer_999 <= lineBuffer_998;
    end
    if (sel) begin
      lineBuffer_1000 <= lineBuffer_999;
    end
    if (sel) begin
      lineBuffer_1001 <= lineBuffer_1000;
    end
    if (sel) begin
      lineBuffer_1002 <= lineBuffer_1001;
    end
    if (sel) begin
      lineBuffer_1003 <= lineBuffer_1002;
    end
    if (sel) begin
      lineBuffer_1004 <= lineBuffer_1003;
    end
    if (sel) begin
      lineBuffer_1005 <= lineBuffer_1004;
    end
    if (sel) begin
      lineBuffer_1006 <= lineBuffer_1005;
    end
    if (sel) begin
      lineBuffer_1007 <= lineBuffer_1006;
    end
    if (sel) begin
      lineBuffer_1008 <= lineBuffer_1007;
    end
    if (sel) begin
      lineBuffer_1009 <= lineBuffer_1008;
    end
    if (sel) begin
      lineBuffer_1010 <= lineBuffer_1009;
    end
    if (sel) begin
      lineBuffer_1011 <= lineBuffer_1010;
    end
    if (sel) begin
      lineBuffer_1012 <= lineBuffer_1011;
    end
    if (sel) begin
      lineBuffer_1013 <= lineBuffer_1012;
    end
    if (sel) begin
      lineBuffer_1014 <= lineBuffer_1013;
    end
    if (sel) begin
      lineBuffer_1015 <= lineBuffer_1014;
    end
    if (sel) begin
      lineBuffer_1016 <= lineBuffer_1015;
    end
    if (sel) begin
      lineBuffer_1017 <= lineBuffer_1016;
    end
    if (sel) begin
      lineBuffer_1018 <= lineBuffer_1017;
    end
    if (sel) begin
      lineBuffer_1019 <= lineBuffer_1018;
    end
    if (sel) begin
      lineBuffer_1020 <= lineBuffer_1019;
    end
    if (sel) begin
      lineBuffer_1021 <= lineBuffer_1020;
    end
    if (sel) begin
      lineBuffer_1022 <= lineBuffer_1021;
    end
    if (sel) begin
      lineBuffer_1023 <= lineBuffer_1022;
    end
    if (sel) begin
      lineBuffer_1024 <= lineBuffer_1023;
    end
    if (sel) begin
      lineBuffer_1025 <= lineBuffer_1024;
    end
    if (sel) begin
      lineBuffer_1026 <= lineBuffer_1025;
    end
    if (sel) begin
      lineBuffer_1027 <= lineBuffer_1026;
    end
    if (sel) begin
      lineBuffer_1028 <= lineBuffer_1027;
    end
    if (sel) begin
      lineBuffer_1029 <= lineBuffer_1028;
    end
    if (sel) begin
      lineBuffer_1030 <= lineBuffer_1029;
    end
    if (sel) begin
      lineBuffer_1031 <= lineBuffer_1030;
    end
    if (sel) begin
      lineBuffer_1032 <= lineBuffer_1031;
    end
    if (sel) begin
      lineBuffer_1033 <= lineBuffer_1032;
    end
    if (sel) begin
      lineBuffer_1034 <= lineBuffer_1033;
    end
    if (sel) begin
      lineBuffer_1035 <= lineBuffer_1034;
    end
    if (sel) begin
      lineBuffer_1036 <= lineBuffer_1035;
    end
    if (sel) begin
      lineBuffer_1037 <= lineBuffer_1036;
    end
    if (sel) begin
      lineBuffer_1038 <= lineBuffer_1037;
    end
    if (sel) begin
      lineBuffer_1039 <= lineBuffer_1038;
    end
    if (sel) begin
      lineBuffer_1040 <= lineBuffer_1039;
    end
    if (sel) begin
      lineBuffer_1041 <= lineBuffer_1040;
    end
    if (sel) begin
      lineBuffer_1042 <= lineBuffer_1041;
    end
    if (sel) begin
      lineBuffer_1043 <= lineBuffer_1042;
    end
    if (sel) begin
      lineBuffer_1044 <= lineBuffer_1043;
    end
    if (sel) begin
      lineBuffer_1045 <= lineBuffer_1044;
    end
    if (sel) begin
      lineBuffer_1046 <= lineBuffer_1045;
    end
    if (sel) begin
      lineBuffer_1047 <= lineBuffer_1046;
    end
    if (sel) begin
      lineBuffer_1048 <= lineBuffer_1047;
    end
    if (sel) begin
      lineBuffer_1049 <= lineBuffer_1048;
    end
    if (sel) begin
      lineBuffer_1050 <= lineBuffer_1049;
    end
    if (sel) begin
      lineBuffer_1051 <= lineBuffer_1050;
    end
    if (sel) begin
      lineBuffer_1052 <= lineBuffer_1051;
    end
    if (sel) begin
      lineBuffer_1053 <= lineBuffer_1052;
    end
    if (sel) begin
      lineBuffer_1054 <= lineBuffer_1053;
    end
    if (sel) begin
      lineBuffer_1055 <= lineBuffer_1054;
    end
    if (sel) begin
      lineBuffer_1056 <= lineBuffer_1055;
    end
    if (sel) begin
      lineBuffer_1057 <= lineBuffer_1056;
    end
    if (sel) begin
      lineBuffer_1058 <= lineBuffer_1057;
    end
    if (sel) begin
      lineBuffer_1059 <= lineBuffer_1058;
    end
    if (sel) begin
      lineBuffer_1060 <= lineBuffer_1059;
    end
    if (sel) begin
      lineBuffer_1061 <= lineBuffer_1060;
    end
    if (sel) begin
      lineBuffer_1062 <= lineBuffer_1061;
    end
    if (sel) begin
      lineBuffer_1063 <= lineBuffer_1062;
    end
    if (sel) begin
      lineBuffer_1064 <= lineBuffer_1063;
    end
    if (sel) begin
      lineBuffer_1065 <= lineBuffer_1064;
    end
    if (sel) begin
      lineBuffer_1066 <= lineBuffer_1065;
    end
    if (sel) begin
      lineBuffer_1067 <= lineBuffer_1066;
    end
    if (sel) begin
      lineBuffer_1068 <= lineBuffer_1067;
    end
    if (sel) begin
      lineBuffer_1069 <= lineBuffer_1068;
    end
    if (sel) begin
      lineBuffer_1070 <= lineBuffer_1069;
    end
    if (sel) begin
      lineBuffer_1071 <= lineBuffer_1070;
    end
    if (sel) begin
      lineBuffer_1072 <= lineBuffer_1071;
    end
    if (sel) begin
      lineBuffer_1073 <= lineBuffer_1072;
    end
    if (sel) begin
      lineBuffer_1074 <= lineBuffer_1073;
    end
    if (sel) begin
      lineBuffer_1075 <= lineBuffer_1074;
    end
    if (sel) begin
      lineBuffer_1076 <= lineBuffer_1075;
    end
    if (sel) begin
      lineBuffer_1077 <= lineBuffer_1076;
    end
    if (sel) begin
      lineBuffer_1078 <= lineBuffer_1077;
    end
    if (sel) begin
      lineBuffer_1079 <= lineBuffer_1078;
    end
    if (sel) begin
      lineBuffer_1080 <= lineBuffer_1079;
    end
    if (sel) begin
      lineBuffer_1081 <= lineBuffer_1080;
    end
    if (sel) begin
      lineBuffer_1082 <= lineBuffer_1081;
    end
    if (sel) begin
      lineBuffer_1083 <= lineBuffer_1082;
    end
    if (sel) begin
      lineBuffer_1084 <= lineBuffer_1083;
    end
    if (sel) begin
      lineBuffer_1085 <= lineBuffer_1084;
    end
    if (sel) begin
      lineBuffer_1086 <= lineBuffer_1085;
    end
    if (sel) begin
      lineBuffer_1087 <= lineBuffer_1086;
    end
    if (sel) begin
      lineBuffer_1088 <= lineBuffer_1087;
    end
    if (sel) begin
      lineBuffer_1089 <= lineBuffer_1088;
    end
    if (sel) begin
      lineBuffer_1090 <= lineBuffer_1089;
    end
    if (sel) begin
      lineBuffer_1091 <= lineBuffer_1090;
    end
    if (sel) begin
      lineBuffer_1092 <= lineBuffer_1091;
    end
    if (sel) begin
      lineBuffer_1093 <= lineBuffer_1092;
    end
    if (sel) begin
      lineBuffer_1094 <= lineBuffer_1093;
    end
    if (sel) begin
      lineBuffer_1095 <= lineBuffer_1094;
    end
    if (sel) begin
      lineBuffer_1096 <= lineBuffer_1095;
    end
    if (sel) begin
      lineBuffer_1097 <= lineBuffer_1096;
    end
    if (sel) begin
      lineBuffer_1098 <= lineBuffer_1097;
    end
    if (sel) begin
      lineBuffer_1099 <= lineBuffer_1098;
    end
    if (sel) begin
      lineBuffer_1100 <= lineBuffer_1099;
    end
    if (sel) begin
      lineBuffer_1101 <= lineBuffer_1100;
    end
    if (sel) begin
      lineBuffer_1102 <= lineBuffer_1101;
    end
    if (sel) begin
      lineBuffer_1103 <= lineBuffer_1102;
    end
    if (sel) begin
      lineBuffer_1104 <= lineBuffer_1103;
    end
    if (sel) begin
      lineBuffer_1105 <= lineBuffer_1104;
    end
    if (sel) begin
      lineBuffer_1106 <= lineBuffer_1105;
    end
    if (sel) begin
      lineBuffer_1107 <= lineBuffer_1106;
    end
    if (sel) begin
      lineBuffer_1108 <= lineBuffer_1107;
    end
    if (sel) begin
      lineBuffer_1109 <= lineBuffer_1108;
    end
    if (sel) begin
      lineBuffer_1110 <= lineBuffer_1109;
    end
    if (sel) begin
      lineBuffer_1111 <= lineBuffer_1110;
    end
    if (sel) begin
      lineBuffer_1112 <= lineBuffer_1111;
    end
    if (sel) begin
      lineBuffer_1113 <= lineBuffer_1112;
    end
    if (sel) begin
      lineBuffer_1114 <= lineBuffer_1113;
    end
    if (sel) begin
      lineBuffer_1115 <= lineBuffer_1114;
    end
    if (sel) begin
      lineBuffer_1116 <= lineBuffer_1115;
    end
    if (sel) begin
      lineBuffer_1117 <= lineBuffer_1116;
    end
    if (sel) begin
      lineBuffer_1118 <= lineBuffer_1117;
    end
    if (sel) begin
      lineBuffer_1119 <= lineBuffer_1118;
    end
    if (sel) begin
      lineBuffer_1120 <= lineBuffer_1119;
    end
    if (sel) begin
      lineBuffer_1121 <= lineBuffer_1120;
    end
    if (sel) begin
      lineBuffer_1122 <= lineBuffer_1121;
    end
    if (sel) begin
      lineBuffer_1123 <= lineBuffer_1122;
    end
    if (sel) begin
      lineBuffer_1124 <= lineBuffer_1123;
    end
    if (sel) begin
      lineBuffer_1125 <= lineBuffer_1124;
    end
    if (sel) begin
      lineBuffer_1126 <= lineBuffer_1125;
    end
    if (sel) begin
      lineBuffer_1127 <= lineBuffer_1126;
    end
    if (sel) begin
      lineBuffer_1128 <= lineBuffer_1127;
    end
    if (sel) begin
      lineBuffer_1129 <= lineBuffer_1128;
    end
    if (sel) begin
      lineBuffer_1130 <= lineBuffer_1129;
    end
    if (sel) begin
      lineBuffer_1131 <= lineBuffer_1130;
    end
    if (sel) begin
      lineBuffer_1132 <= lineBuffer_1131;
    end
    if (sel) begin
      lineBuffer_1133 <= lineBuffer_1132;
    end
    if (sel) begin
      lineBuffer_1134 <= lineBuffer_1133;
    end
    if (sel) begin
      lineBuffer_1135 <= lineBuffer_1134;
    end
    if (sel) begin
      lineBuffer_1136 <= lineBuffer_1135;
    end
    if (sel) begin
      lineBuffer_1137 <= lineBuffer_1136;
    end
    if (sel) begin
      lineBuffer_1138 <= lineBuffer_1137;
    end
    if (sel) begin
      lineBuffer_1139 <= lineBuffer_1138;
    end
    if (sel) begin
      lineBuffer_1140 <= lineBuffer_1139;
    end
    if (sel) begin
      lineBuffer_1141 <= lineBuffer_1140;
    end
    if (sel) begin
      lineBuffer_1142 <= lineBuffer_1141;
    end
    if (sel) begin
      lineBuffer_1143 <= lineBuffer_1142;
    end
    if (sel) begin
      lineBuffer_1144 <= lineBuffer_1143;
    end
    if (sel) begin
      lineBuffer_1145 <= lineBuffer_1144;
    end
    if (sel) begin
      lineBuffer_1146 <= lineBuffer_1145;
    end
    if (sel) begin
      lineBuffer_1147 <= lineBuffer_1146;
    end
    if (sel) begin
      lineBuffer_1148 <= lineBuffer_1147;
    end
    if (sel) begin
      lineBuffer_1149 <= lineBuffer_1148;
    end
    if (sel) begin
      lineBuffer_1150 <= lineBuffer_1149;
    end
    if (sel) begin
      lineBuffer_1151 <= lineBuffer_1150;
    end
    if (sel) begin
      lineBuffer_1152 <= lineBuffer_1151;
    end
    if (sel) begin
      lineBuffer_1153 <= lineBuffer_1152;
    end
    if (sel) begin
      lineBuffer_1154 <= lineBuffer_1153;
    end
    if (sel) begin
      lineBuffer_1155 <= lineBuffer_1154;
    end
    if (sel) begin
      lineBuffer_1156 <= lineBuffer_1155;
    end
    if (sel) begin
      lineBuffer_1157 <= lineBuffer_1156;
    end
    if (sel) begin
      lineBuffer_1158 <= lineBuffer_1157;
    end
    if (sel) begin
      lineBuffer_1159 <= lineBuffer_1158;
    end
    if (sel) begin
      lineBuffer_1160 <= lineBuffer_1159;
    end
    if (sel) begin
      lineBuffer_1161 <= lineBuffer_1160;
    end
    if (sel) begin
      lineBuffer_1162 <= lineBuffer_1161;
    end
    if (sel) begin
      lineBuffer_1163 <= lineBuffer_1162;
    end
    if (sel) begin
      lineBuffer_1164 <= lineBuffer_1163;
    end
    if (sel) begin
      lineBuffer_1165 <= lineBuffer_1164;
    end
    if (sel) begin
      lineBuffer_1166 <= lineBuffer_1165;
    end
    if (sel) begin
      lineBuffer_1167 <= lineBuffer_1166;
    end
    if (sel) begin
      lineBuffer_1168 <= lineBuffer_1167;
    end
    if (sel) begin
      lineBuffer_1169 <= lineBuffer_1168;
    end
    if (sel) begin
      lineBuffer_1170 <= lineBuffer_1169;
    end
    if (sel) begin
      lineBuffer_1171 <= lineBuffer_1170;
    end
    if (sel) begin
      lineBuffer_1172 <= lineBuffer_1171;
    end
    if (sel) begin
      lineBuffer_1173 <= lineBuffer_1172;
    end
    if (sel) begin
      lineBuffer_1174 <= lineBuffer_1173;
    end
    if (sel) begin
      lineBuffer_1175 <= lineBuffer_1174;
    end
    if (sel) begin
      lineBuffer_1176 <= lineBuffer_1175;
    end
    if (sel) begin
      lineBuffer_1177 <= lineBuffer_1176;
    end
    if (sel) begin
      lineBuffer_1178 <= lineBuffer_1177;
    end
    if (sel) begin
      lineBuffer_1179 <= lineBuffer_1178;
    end
    if (sel) begin
      lineBuffer_1180 <= lineBuffer_1179;
    end
    if (sel) begin
      lineBuffer_1181 <= lineBuffer_1180;
    end
    if (sel) begin
      lineBuffer_1182 <= lineBuffer_1181;
    end
    if (sel) begin
      lineBuffer_1183 <= lineBuffer_1182;
    end
    if (sel) begin
      lineBuffer_1184 <= lineBuffer_1183;
    end
    if (sel) begin
      lineBuffer_1185 <= lineBuffer_1184;
    end
    if (sel) begin
      lineBuffer_1186 <= lineBuffer_1185;
    end
    if (sel) begin
      lineBuffer_1187 <= lineBuffer_1186;
    end
    if (sel) begin
      lineBuffer_1188 <= lineBuffer_1187;
    end
    if (sel) begin
      lineBuffer_1189 <= lineBuffer_1188;
    end
    if (sel) begin
      lineBuffer_1190 <= lineBuffer_1189;
    end
    if (sel) begin
      lineBuffer_1191 <= lineBuffer_1190;
    end
    if (sel) begin
      lineBuffer_1192 <= lineBuffer_1191;
    end
    if (sel) begin
      lineBuffer_1193 <= lineBuffer_1192;
    end
    if (sel) begin
      lineBuffer_1194 <= lineBuffer_1193;
    end
    if (sel) begin
      lineBuffer_1195 <= lineBuffer_1194;
    end
    if (sel) begin
      lineBuffer_1196 <= lineBuffer_1195;
    end
    if (sel) begin
      lineBuffer_1197 <= lineBuffer_1196;
    end
    if (sel) begin
      lineBuffer_1198 <= lineBuffer_1197;
    end
    if (sel) begin
      lineBuffer_1199 <= lineBuffer_1198;
    end
    if (sel) begin
      lineBuffer_1200 <= lineBuffer_1199;
    end
    if (sel) begin
      lineBuffer_1201 <= lineBuffer_1200;
    end
    if (sel) begin
      lineBuffer_1202 <= lineBuffer_1201;
    end
    if (sel) begin
      lineBuffer_1203 <= lineBuffer_1202;
    end
    if (sel) begin
      lineBuffer_1204 <= lineBuffer_1203;
    end
    if (sel) begin
      lineBuffer_1205 <= lineBuffer_1204;
    end
    if (sel) begin
      lineBuffer_1206 <= lineBuffer_1205;
    end
    if (sel) begin
      lineBuffer_1207 <= lineBuffer_1206;
    end
    if (sel) begin
      lineBuffer_1208 <= lineBuffer_1207;
    end
    if (sel) begin
      lineBuffer_1209 <= lineBuffer_1208;
    end
    if (sel) begin
      lineBuffer_1210 <= lineBuffer_1209;
    end
    if (sel) begin
      lineBuffer_1211 <= lineBuffer_1210;
    end
    if (sel) begin
      lineBuffer_1212 <= lineBuffer_1211;
    end
    if (sel) begin
      lineBuffer_1213 <= lineBuffer_1212;
    end
    if (sel) begin
      lineBuffer_1214 <= lineBuffer_1213;
    end
    if (sel) begin
      lineBuffer_1215 <= lineBuffer_1214;
    end
    if (sel) begin
      lineBuffer_1216 <= lineBuffer_1215;
    end
    if (sel) begin
      lineBuffer_1217 <= lineBuffer_1216;
    end
    if (sel) begin
      lineBuffer_1218 <= lineBuffer_1217;
    end
    if (sel) begin
      lineBuffer_1219 <= lineBuffer_1218;
    end
    if (sel) begin
      lineBuffer_1220 <= lineBuffer_1219;
    end
    if (sel) begin
      lineBuffer_1221 <= lineBuffer_1220;
    end
    if (sel) begin
      lineBuffer_1222 <= lineBuffer_1221;
    end
    if (sel) begin
      lineBuffer_1223 <= lineBuffer_1222;
    end
    if (sel) begin
      lineBuffer_1224 <= lineBuffer_1223;
    end
    if (sel) begin
      lineBuffer_1225 <= lineBuffer_1224;
    end
    if (sel) begin
      lineBuffer_1226 <= lineBuffer_1225;
    end
    if (sel) begin
      lineBuffer_1227 <= lineBuffer_1226;
    end
    if (sel) begin
      lineBuffer_1228 <= lineBuffer_1227;
    end
    if (sel) begin
      lineBuffer_1229 <= lineBuffer_1228;
    end
    if (sel) begin
      lineBuffer_1230 <= lineBuffer_1229;
    end
    if (sel) begin
      lineBuffer_1231 <= lineBuffer_1230;
    end
    if (sel) begin
      lineBuffer_1232 <= lineBuffer_1231;
    end
    if (sel) begin
      lineBuffer_1233 <= lineBuffer_1232;
    end
    if (sel) begin
      lineBuffer_1234 <= lineBuffer_1233;
    end
    if (sel) begin
      lineBuffer_1235 <= lineBuffer_1234;
    end
    if (sel) begin
      lineBuffer_1236 <= lineBuffer_1235;
    end
    if (sel) begin
      lineBuffer_1237 <= lineBuffer_1236;
    end
    if (sel) begin
      lineBuffer_1238 <= lineBuffer_1237;
    end
    if (sel) begin
      lineBuffer_1239 <= lineBuffer_1238;
    end
    if (sel) begin
      lineBuffer_1240 <= lineBuffer_1239;
    end
    if (sel) begin
      lineBuffer_1241 <= lineBuffer_1240;
    end
    if (sel) begin
      lineBuffer_1242 <= lineBuffer_1241;
    end
    if (sel) begin
      lineBuffer_1243 <= lineBuffer_1242;
    end
    if (sel) begin
      lineBuffer_1244 <= lineBuffer_1243;
    end
    if (sel) begin
      lineBuffer_1245 <= lineBuffer_1244;
    end
    if (sel) begin
      lineBuffer_1246 <= lineBuffer_1245;
    end
    if (sel) begin
      lineBuffer_1247 <= lineBuffer_1246;
    end
    if (sel) begin
      lineBuffer_1248 <= lineBuffer_1247;
    end
    if (sel) begin
      lineBuffer_1249 <= lineBuffer_1248;
    end
    if (sel) begin
      lineBuffer_1250 <= lineBuffer_1249;
    end
    if (sel) begin
      lineBuffer_1251 <= lineBuffer_1250;
    end
    if (sel) begin
      lineBuffer_1252 <= lineBuffer_1251;
    end
    if (sel) begin
      lineBuffer_1253 <= lineBuffer_1252;
    end
    if (sel) begin
      lineBuffer_1254 <= lineBuffer_1253;
    end
    if (sel) begin
      lineBuffer_1255 <= lineBuffer_1254;
    end
    if (sel) begin
      lineBuffer_1256 <= lineBuffer_1255;
    end
    if (sel) begin
      lineBuffer_1257 <= lineBuffer_1256;
    end
    if (sel) begin
      lineBuffer_1258 <= lineBuffer_1257;
    end
    if (sel) begin
      lineBuffer_1259 <= lineBuffer_1258;
    end
    if (sel) begin
      lineBuffer_1260 <= lineBuffer_1259;
    end
    if (sel) begin
      lineBuffer_1261 <= lineBuffer_1260;
    end
    if (sel) begin
      lineBuffer_1262 <= lineBuffer_1261;
    end
    if (sel) begin
      lineBuffer_1263 <= lineBuffer_1262;
    end
    if (sel) begin
      lineBuffer_1264 <= lineBuffer_1263;
    end
    if (sel) begin
      lineBuffer_1265 <= lineBuffer_1264;
    end
    if (sel) begin
      lineBuffer_1266 <= lineBuffer_1265;
    end
    if (sel) begin
      lineBuffer_1267 <= lineBuffer_1266;
    end
    if (sel) begin
      lineBuffer_1268 <= lineBuffer_1267;
    end
    if (sel) begin
      lineBuffer_1269 <= lineBuffer_1268;
    end
    if (sel) begin
      lineBuffer_1270 <= lineBuffer_1269;
    end
    if (sel) begin
      lineBuffer_1271 <= lineBuffer_1270;
    end
    if (sel) begin
      lineBuffer_1272 <= lineBuffer_1271;
    end
    if (sel) begin
      lineBuffer_1273 <= lineBuffer_1272;
    end
    if (sel) begin
      lineBuffer_1274 <= lineBuffer_1273;
    end
    if (sel) begin
      lineBuffer_1275 <= lineBuffer_1274;
    end
    if (sel) begin
      lineBuffer_1276 <= lineBuffer_1275;
    end
    if (sel) begin
      lineBuffer_1277 <= lineBuffer_1276;
    end
    if (sel) begin
      lineBuffer_1278 <= lineBuffer_1277;
    end
    if (sel) begin
      lineBuffer_1279 <= lineBuffer_1278;
    end
    if (sel) begin
      lineBuffer_1280 <= lineBuffer_1279;
    end
    if (sel) begin
      lineBuffer_1281 <= lineBuffer_1280;
    end
    if (sel) begin
      lineBuffer_1282 <= lineBuffer_1281;
    end
    if (sel) begin
      lineBuffer_1283 <= lineBuffer_1282;
    end
    if (sel) begin
      lineBuffer_1284 <= lineBuffer_1283;
    end
    if (sel) begin
      lineBuffer_1285 <= lineBuffer_1284;
    end
    if (sel) begin
      lineBuffer_1286 <= lineBuffer_1285;
    end
    if (sel) begin
      lineBuffer_1287 <= lineBuffer_1286;
    end
    if (sel) begin
      lineBuffer_1288 <= lineBuffer_1287;
    end
    if (sel) begin
      lineBuffer_1289 <= lineBuffer_1288;
    end
    if (sel) begin
      lineBuffer_1290 <= lineBuffer_1289;
    end
    if (sel) begin
      lineBuffer_1291 <= lineBuffer_1290;
    end
    if (sel) begin
      lineBuffer_1292 <= lineBuffer_1291;
    end
    if (sel) begin
      lineBuffer_1293 <= lineBuffer_1292;
    end
    if (sel) begin
      lineBuffer_1294 <= lineBuffer_1293;
    end
    if (sel) begin
      lineBuffer_1295 <= lineBuffer_1294;
    end
    if (sel) begin
      lineBuffer_1296 <= lineBuffer_1295;
    end
    if (sel) begin
      lineBuffer_1297 <= lineBuffer_1296;
    end
    if (sel) begin
      lineBuffer_1298 <= lineBuffer_1297;
    end
    if (sel) begin
      lineBuffer_1299 <= lineBuffer_1298;
    end
    if (sel) begin
      lineBuffer_1300 <= lineBuffer_1299;
    end
    if (sel) begin
      lineBuffer_1301 <= lineBuffer_1300;
    end
    if (sel) begin
      lineBuffer_1302 <= lineBuffer_1301;
    end
    if (sel) begin
      lineBuffer_1303 <= lineBuffer_1302;
    end
    if (sel) begin
      lineBuffer_1304 <= lineBuffer_1303;
    end
    if (sel) begin
      lineBuffer_1305 <= lineBuffer_1304;
    end
    if (sel) begin
      lineBuffer_1306 <= lineBuffer_1305;
    end
    if (sel) begin
      lineBuffer_1307 <= lineBuffer_1306;
    end
    if (sel) begin
      lineBuffer_1308 <= lineBuffer_1307;
    end
    if (sel) begin
      lineBuffer_1309 <= lineBuffer_1308;
    end
    if (sel) begin
      lineBuffer_1310 <= lineBuffer_1309;
    end
    if (sel) begin
      lineBuffer_1311 <= lineBuffer_1310;
    end
    if (sel) begin
      lineBuffer_1312 <= lineBuffer_1311;
    end
    if (sel) begin
      lineBuffer_1313 <= lineBuffer_1312;
    end
    if (sel) begin
      lineBuffer_1314 <= lineBuffer_1313;
    end
    if (sel) begin
      lineBuffer_1315 <= lineBuffer_1314;
    end
    if (sel) begin
      lineBuffer_1316 <= lineBuffer_1315;
    end
    if (sel) begin
      lineBuffer_1317 <= lineBuffer_1316;
    end
    if (sel) begin
      lineBuffer_1318 <= lineBuffer_1317;
    end
    if (sel) begin
      lineBuffer_1319 <= lineBuffer_1318;
    end
    if (sel) begin
      lineBuffer_1320 <= lineBuffer_1319;
    end
    if (sel) begin
      lineBuffer_1321 <= lineBuffer_1320;
    end
    if (sel) begin
      lineBuffer_1322 <= lineBuffer_1321;
    end
    if (sel) begin
      lineBuffer_1323 <= lineBuffer_1322;
    end
    if (sel) begin
      lineBuffer_1324 <= lineBuffer_1323;
    end
    if (sel) begin
      lineBuffer_1325 <= lineBuffer_1324;
    end
    if (sel) begin
      lineBuffer_1326 <= lineBuffer_1325;
    end
    if (sel) begin
      lineBuffer_1327 <= lineBuffer_1326;
    end
    if (sel) begin
      lineBuffer_1328 <= lineBuffer_1327;
    end
    if (sel) begin
      lineBuffer_1329 <= lineBuffer_1328;
    end
    if (sel) begin
      lineBuffer_1330 <= lineBuffer_1329;
    end
    if (sel) begin
      lineBuffer_1331 <= lineBuffer_1330;
    end
    if (sel) begin
      lineBuffer_1332 <= lineBuffer_1331;
    end
    if (sel) begin
      lineBuffer_1333 <= lineBuffer_1332;
    end
    if (sel) begin
      lineBuffer_1334 <= lineBuffer_1333;
    end
    if (sel) begin
      lineBuffer_1335 <= lineBuffer_1334;
    end
    if (sel) begin
      lineBuffer_1336 <= lineBuffer_1335;
    end
    if (sel) begin
      lineBuffer_1337 <= lineBuffer_1336;
    end
    if (sel) begin
      lineBuffer_1338 <= lineBuffer_1337;
    end
    if (sel) begin
      lineBuffer_1339 <= lineBuffer_1338;
    end
    if (sel) begin
      lineBuffer_1340 <= lineBuffer_1339;
    end
    if (sel) begin
      lineBuffer_1341 <= lineBuffer_1340;
    end
    if (sel) begin
      lineBuffer_1342 <= lineBuffer_1341;
    end
    if (sel) begin
      lineBuffer_1343 <= lineBuffer_1342;
    end
    if (sel) begin
      lineBuffer_1344 <= lineBuffer_1343;
    end
    if (sel) begin
      lineBuffer_1345 <= lineBuffer_1344;
    end
    if (sel) begin
      lineBuffer_1346 <= lineBuffer_1345;
    end
    if (sel) begin
      lineBuffer_1347 <= lineBuffer_1346;
    end
    if (sel) begin
      lineBuffer_1348 <= lineBuffer_1347;
    end
    if (sel) begin
      lineBuffer_1349 <= lineBuffer_1348;
    end
    if (sel) begin
      lineBuffer_1350 <= lineBuffer_1349;
    end
    if (sel) begin
      lineBuffer_1351 <= lineBuffer_1350;
    end
    if (sel) begin
      lineBuffer_1352 <= lineBuffer_1351;
    end
    if (sel) begin
      lineBuffer_1353 <= lineBuffer_1352;
    end
    if (sel) begin
      lineBuffer_1354 <= lineBuffer_1353;
    end
    if (sel) begin
      lineBuffer_1355 <= lineBuffer_1354;
    end
    if (sel) begin
      lineBuffer_1356 <= lineBuffer_1355;
    end
    if (sel) begin
      lineBuffer_1357 <= lineBuffer_1356;
    end
    if (sel) begin
      lineBuffer_1358 <= lineBuffer_1357;
    end
    if (sel) begin
      lineBuffer_1359 <= lineBuffer_1358;
    end
    if (sel) begin
      lineBuffer_1360 <= lineBuffer_1359;
    end
    if (sel) begin
      lineBuffer_1361 <= lineBuffer_1360;
    end
    if (sel) begin
      lineBuffer_1362 <= lineBuffer_1361;
    end
    if (sel) begin
      lineBuffer_1363 <= lineBuffer_1362;
    end
    if (sel) begin
      lineBuffer_1364 <= lineBuffer_1363;
    end
    if (sel) begin
      lineBuffer_1365 <= lineBuffer_1364;
    end
    if (sel) begin
      lineBuffer_1366 <= lineBuffer_1365;
    end
    if (sel) begin
      lineBuffer_1367 <= lineBuffer_1366;
    end
    if (sel) begin
      lineBuffer_1368 <= lineBuffer_1367;
    end
    if (sel) begin
      lineBuffer_1369 <= lineBuffer_1368;
    end
    if (sel) begin
      lineBuffer_1370 <= lineBuffer_1369;
    end
    if (sel) begin
      lineBuffer_1371 <= lineBuffer_1370;
    end
    if (sel) begin
      lineBuffer_1372 <= lineBuffer_1371;
    end
    if (sel) begin
      lineBuffer_1373 <= lineBuffer_1372;
    end
    if (sel) begin
      lineBuffer_1374 <= lineBuffer_1373;
    end
    if (sel) begin
      lineBuffer_1375 <= lineBuffer_1374;
    end
    if (sel) begin
      lineBuffer_1376 <= lineBuffer_1375;
    end
    if (sel) begin
      lineBuffer_1377 <= lineBuffer_1376;
    end
    if (sel) begin
      lineBuffer_1378 <= lineBuffer_1377;
    end
    if (sel) begin
      lineBuffer_1379 <= lineBuffer_1378;
    end
    if (sel) begin
      lineBuffer_1380 <= lineBuffer_1379;
    end
    if (sel) begin
      lineBuffer_1381 <= lineBuffer_1380;
    end
    if (sel) begin
      lineBuffer_1382 <= lineBuffer_1381;
    end
    if (sel) begin
      lineBuffer_1383 <= lineBuffer_1382;
    end
    if (sel) begin
      lineBuffer_1384 <= lineBuffer_1383;
    end
    if (sel) begin
      lineBuffer_1385 <= lineBuffer_1384;
    end
    if (sel) begin
      lineBuffer_1386 <= lineBuffer_1385;
    end
    if (sel) begin
      lineBuffer_1387 <= lineBuffer_1386;
    end
    if (sel) begin
      lineBuffer_1388 <= lineBuffer_1387;
    end
    if (sel) begin
      lineBuffer_1389 <= lineBuffer_1388;
    end
    if (sel) begin
      lineBuffer_1390 <= lineBuffer_1389;
    end
    if (sel) begin
      lineBuffer_1391 <= lineBuffer_1390;
    end
    if (sel) begin
      lineBuffer_1392 <= lineBuffer_1391;
    end
    if (sel) begin
      lineBuffer_1393 <= lineBuffer_1392;
    end
    if (sel) begin
      lineBuffer_1394 <= lineBuffer_1393;
    end
    if (sel) begin
      lineBuffer_1395 <= lineBuffer_1394;
    end
    if (sel) begin
      lineBuffer_1396 <= lineBuffer_1395;
    end
    if (sel) begin
      lineBuffer_1397 <= lineBuffer_1396;
    end
    if (sel) begin
      lineBuffer_1398 <= lineBuffer_1397;
    end
    if (sel) begin
      lineBuffer_1399 <= lineBuffer_1398;
    end
    if (sel) begin
      lineBuffer_1400 <= lineBuffer_1399;
    end
    if (sel) begin
      lineBuffer_1401 <= lineBuffer_1400;
    end
    if (sel) begin
      lineBuffer_1402 <= lineBuffer_1401;
    end
    if (sel) begin
      lineBuffer_1403 <= lineBuffer_1402;
    end
    if (sel) begin
      lineBuffer_1404 <= lineBuffer_1403;
    end
    if (sel) begin
      lineBuffer_1405 <= lineBuffer_1404;
    end
    if (sel) begin
      lineBuffer_1406 <= lineBuffer_1405;
    end
    if (sel) begin
      lineBuffer_1407 <= lineBuffer_1406;
    end
    if (sel) begin
      lineBuffer_1408 <= lineBuffer_1407;
    end
    if (sel) begin
      lineBuffer_1409 <= lineBuffer_1408;
    end
    if (sel) begin
      lineBuffer_1410 <= lineBuffer_1409;
    end
    if (sel) begin
      lineBuffer_1411 <= lineBuffer_1410;
    end
    if (sel) begin
      lineBuffer_1412 <= lineBuffer_1411;
    end
    if (sel) begin
      lineBuffer_1413 <= lineBuffer_1412;
    end
    if (sel) begin
      lineBuffer_1414 <= lineBuffer_1413;
    end
    if (sel) begin
      lineBuffer_1415 <= lineBuffer_1414;
    end
    if (sel) begin
      lineBuffer_1416 <= lineBuffer_1415;
    end
    if (sel) begin
      lineBuffer_1417 <= lineBuffer_1416;
    end
    if (sel) begin
      lineBuffer_1418 <= lineBuffer_1417;
    end
    if (sel) begin
      lineBuffer_1419 <= lineBuffer_1418;
    end
    if (sel) begin
      lineBuffer_1420 <= lineBuffer_1419;
    end
    if (sel) begin
      lineBuffer_1421 <= lineBuffer_1420;
    end
    if (sel) begin
      lineBuffer_1422 <= lineBuffer_1421;
    end
    if (sel) begin
      lineBuffer_1423 <= lineBuffer_1422;
    end
    if (sel) begin
      lineBuffer_1424 <= lineBuffer_1423;
    end
    if (sel) begin
      lineBuffer_1425 <= lineBuffer_1424;
    end
    if (sel) begin
      lineBuffer_1426 <= lineBuffer_1425;
    end
    if (sel) begin
      lineBuffer_1427 <= lineBuffer_1426;
    end
    if (sel) begin
      lineBuffer_1428 <= lineBuffer_1427;
    end
    if (sel) begin
      lineBuffer_1429 <= lineBuffer_1428;
    end
    if (sel) begin
      lineBuffer_1430 <= lineBuffer_1429;
    end
    if (sel) begin
      lineBuffer_1431 <= lineBuffer_1430;
    end
    if (sel) begin
      lineBuffer_1432 <= lineBuffer_1431;
    end
    if (sel) begin
      lineBuffer_1433 <= lineBuffer_1432;
    end
    if (sel) begin
      lineBuffer_1434 <= lineBuffer_1433;
    end
    if (sel) begin
      lineBuffer_1435 <= lineBuffer_1434;
    end
    if (sel) begin
      lineBuffer_1436 <= lineBuffer_1435;
    end
    if (sel) begin
      lineBuffer_1437 <= lineBuffer_1436;
    end
    if (sel) begin
      lineBuffer_1438 <= lineBuffer_1437;
    end
    if (sel) begin
      lineBuffer_1439 <= lineBuffer_1438;
    end
    if (sel) begin
      lineBuffer_1440 <= lineBuffer_1439;
    end
    if (sel) begin
      lineBuffer_1441 <= lineBuffer_1440;
    end
    if (sel) begin
      lineBuffer_1442 <= lineBuffer_1441;
    end
    if (sel) begin
      lineBuffer_1443 <= lineBuffer_1442;
    end
    if (sel) begin
      lineBuffer_1444 <= lineBuffer_1443;
    end
    if (sel) begin
      lineBuffer_1445 <= lineBuffer_1444;
    end
    if (sel) begin
      lineBuffer_1446 <= lineBuffer_1445;
    end
    if (sel) begin
      lineBuffer_1447 <= lineBuffer_1446;
    end
    if (sel) begin
      lineBuffer_1448 <= lineBuffer_1447;
    end
    if (sel) begin
      lineBuffer_1449 <= lineBuffer_1448;
    end
    if (sel) begin
      lineBuffer_1450 <= lineBuffer_1449;
    end
    if (sel) begin
      lineBuffer_1451 <= lineBuffer_1450;
    end
    if (sel) begin
      lineBuffer_1452 <= lineBuffer_1451;
    end
    if (sel) begin
      lineBuffer_1453 <= lineBuffer_1452;
    end
    if (sel) begin
      lineBuffer_1454 <= lineBuffer_1453;
    end
    if (sel) begin
      lineBuffer_1455 <= lineBuffer_1454;
    end
    if (sel) begin
      lineBuffer_1456 <= lineBuffer_1455;
    end
    if (sel) begin
      lineBuffer_1457 <= lineBuffer_1456;
    end
    if (sel) begin
      lineBuffer_1458 <= lineBuffer_1457;
    end
    if (sel) begin
      lineBuffer_1459 <= lineBuffer_1458;
    end
    if (sel) begin
      lineBuffer_1460 <= lineBuffer_1459;
    end
    if (sel) begin
      lineBuffer_1461 <= lineBuffer_1460;
    end
    if (sel) begin
      lineBuffer_1462 <= lineBuffer_1461;
    end
    if (sel) begin
      lineBuffer_1463 <= lineBuffer_1462;
    end
    if (sel) begin
      lineBuffer_1464 <= lineBuffer_1463;
    end
    if (sel) begin
      lineBuffer_1465 <= lineBuffer_1464;
    end
    if (sel) begin
      lineBuffer_1466 <= lineBuffer_1465;
    end
    if (sel) begin
      lineBuffer_1467 <= lineBuffer_1466;
    end
    if (sel) begin
      lineBuffer_1468 <= lineBuffer_1467;
    end
    if (sel) begin
      lineBuffer_1469 <= lineBuffer_1468;
    end
    if (sel) begin
      lineBuffer_1470 <= lineBuffer_1469;
    end
    if (sel) begin
      lineBuffer_1471 <= lineBuffer_1470;
    end
    if (sel) begin
      lineBuffer_1472 <= lineBuffer_1471;
    end
    if (sel) begin
      lineBuffer_1473 <= lineBuffer_1472;
    end
    if (sel) begin
      lineBuffer_1474 <= lineBuffer_1473;
    end
    if (sel) begin
      lineBuffer_1475 <= lineBuffer_1474;
    end
    if (sel) begin
      lineBuffer_1476 <= lineBuffer_1475;
    end
    if (sel) begin
      lineBuffer_1477 <= lineBuffer_1476;
    end
    if (sel) begin
      lineBuffer_1478 <= lineBuffer_1477;
    end
    if (sel) begin
      lineBuffer_1479 <= lineBuffer_1478;
    end
    if (sel) begin
      lineBuffer_1480 <= lineBuffer_1479;
    end
    if (sel) begin
      lineBuffer_1481 <= lineBuffer_1480;
    end
    if (sel) begin
      lineBuffer_1482 <= lineBuffer_1481;
    end
    if (sel) begin
      lineBuffer_1483 <= lineBuffer_1482;
    end
    if (sel) begin
      lineBuffer_1484 <= lineBuffer_1483;
    end
    if (sel) begin
      lineBuffer_1485 <= lineBuffer_1484;
    end
    if (sel) begin
      lineBuffer_1486 <= lineBuffer_1485;
    end
    if (sel) begin
      lineBuffer_1487 <= lineBuffer_1486;
    end
    if (sel) begin
      lineBuffer_1488 <= lineBuffer_1487;
    end
    if (sel) begin
      lineBuffer_1489 <= lineBuffer_1488;
    end
    if (sel) begin
      lineBuffer_1490 <= lineBuffer_1489;
    end
    if (sel) begin
      lineBuffer_1491 <= lineBuffer_1490;
    end
    if (sel) begin
      lineBuffer_1492 <= lineBuffer_1491;
    end
    if (sel) begin
      lineBuffer_1493 <= lineBuffer_1492;
    end
    if (sel) begin
      lineBuffer_1494 <= lineBuffer_1493;
    end
    if (sel) begin
      lineBuffer_1495 <= lineBuffer_1494;
    end
    if (sel) begin
      lineBuffer_1496 <= lineBuffer_1495;
    end
    if (sel) begin
      lineBuffer_1497 <= lineBuffer_1496;
    end
    if (sel) begin
      lineBuffer_1498 <= lineBuffer_1497;
    end
    if (sel) begin
      lineBuffer_1499 <= lineBuffer_1498;
    end
    if (sel) begin
      lineBuffer_1500 <= lineBuffer_1499;
    end
    if (sel) begin
      lineBuffer_1501 <= lineBuffer_1500;
    end
    if (sel) begin
      lineBuffer_1502 <= lineBuffer_1501;
    end
    if (sel) begin
      lineBuffer_1503 <= lineBuffer_1502;
    end
    if (sel) begin
      lineBuffer_1504 <= lineBuffer_1503;
    end
    if (sel) begin
      lineBuffer_1505 <= lineBuffer_1504;
    end
    if (sel) begin
      lineBuffer_1506 <= lineBuffer_1505;
    end
    if (sel) begin
      lineBuffer_1507 <= lineBuffer_1506;
    end
    if (sel) begin
      lineBuffer_1508 <= lineBuffer_1507;
    end
    if (sel) begin
      lineBuffer_1509 <= lineBuffer_1508;
    end
    if (sel) begin
      lineBuffer_1510 <= lineBuffer_1509;
    end
    if (sel) begin
      lineBuffer_1511 <= lineBuffer_1510;
    end
    if (sel) begin
      lineBuffer_1512 <= lineBuffer_1511;
    end
    if (sel) begin
      lineBuffer_1513 <= lineBuffer_1512;
    end
    if (sel) begin
      lineBuffer_1514 <= lineBuffer_1513;
    end
    if (sel) begin
      lineBuffer_1515 <= lineBuffer_1514;
    end
    if (sel) begin
      lineBuffer_1516 <= lineBuffer_1515;
    end
    if (sel) begin
      lineBuffer_1517 <= lineBuffer_1516;
    end
    if (sel) begin
      lineBuffer_1518 <= lineBuffer_1517;
    end
    if (sel) begin
      lineBuffer_1519 <= lineBuffer_1518;
    end
    if (sel) begin
      lineBuffer_1520 <= lineBuffer_1519;
    end
    if (sel) begin
      lineBuffer_1521 <= lineBuffer_1520;
    end
    if (sel) begin
      lineBuffer_1522 <= lineBuffer_1521;
    end
    if (sel) begin
      lineBuffer_1523 <= lineBuffer_1522;
    end
    if (sel) begin
      lineBuffer_1524 <= lineBuffer_1523;
    end
    if (sel) begin
      lineBuffer_1525 <= lineBuffer_1524;
    end
    if (sel) begin
      lineBuffer_1526 <= lineBuffer_1525;
    end
    if (sel) begin
      lineBuffer_1527 <= lineBuffer_1526;
    end
    if (sel) begin
      lineBuffer_1528 <= lineBuffer_1527;
    end
    if (sel) begin
      lineBuffer_1529 <= lineBuffer_1528;
    end
    if (sel) begin
      lineBuffer_1530 <= lineBuffer_1529;
    end
    if (sel) begin
      lineBuffer_1531 <= lineBuffer_1530;
    end
    if (sel) begin
      lineBuffer_1532 <= lineBuffer_1531;
    end
    if (sel) begin
      lineBuffer_1533 <= lineBuffer_1532;
    end
    if (sel) begin
      lineBuffer_1534 <= lineBuffer_1533;
    end
    if (sel) begin
      lineBuffer_1535 <= lineBuffer_1534;
    end
    if (sel) begin
      lineBuffer_1536 <= lineBuffer_1535;
    end
    if (sel) begin
      lineBuffer_1537 <= lineBuffer_1536;
    end
    if (sel) begin
      lineBuffer_1538 <= lineBuffer_1537;
    end
    if (sel) begin
      lineBuffer_1539 <= lineBuffer_1538;
    end
    if (sel) begin
      lineBuffer_1540 <= lineBuffer_1539;
    end
    if (sel) begin
      lineBuffer_1541 <= lineBuffer_1540;
    end
    if (sel) begin
      lineBuffer_1542 <= lineBuffer_1541;
    end
    if (sel) begin
      lineBuffer_1543 <= lineBuffer_1542;
    end
    if (sel) begin
      lineBuffer_1544 <= lineBuffer_1543;
    end
    if (sel) begin
      lineBuffer_1545 <= lineBuffer_1544;
    end
    if (sel) begin
      lineBuffer_1546 <= lineBuffer_1545;
    end
    if (sel) begin
      lineBuffer_1547 <= lineBuffer_1546;
    end
    if (sel) begin
      lineBuffer_1548 <= lineBuffer_1547;
    end
    if (sel) begin
      lineBuffer_1549 <= lineBuffer_1548;
    end
    if (sel) begin
      lineBuffer_1550 <= lineBuffer_1549;
    end
    if (sel) begin
      lineBuffer_1551 <= lineBuffer_1550;
    end
    if (sel) begin
      lineBuffer_1552 <= lineBuffer_1551;
    end
    if (sel) begin
      lineBuffer_1553 <= lineBuffer_1552;
    end
    if (sel) begin
      lineBuffer_1554 <= lineBuffer_1553;
    end
    if (sel) begin
      lineBuffer_1555 <= lineBuffer_1554;
    end
    if (sel) begin
      lineBuffer_1556 <= lineBuffer_1555;
    end
    if (sel) begin
      lineBuffer_1557 <= lineBuffer_1556;
    end
    if (sel) begin
      lineBuffer_1558 <= lineBuffer_1557;
    end
    if (sel) begin
      lineBuffer_1559 <= lineBuffer_1558;
    end
    if (sel) begin
      lineBuffer_1560 <= lineBuffer_1559;
    end
    if (sel) begin
      lineBuffer_1561 <= lineBuffer_1560;
    end
    if (sel) begin
      lineBuffer_1562 <= lineBuffer_1561;
    end
    if (sel) begin
      lineBuffer_1563 <= lineBuffer_1562;
    end
    if (sel) begin
      lineBuffer_1564 <= lineBuffer_1563;
    end
    if (sel) begin
      lineBuffer_1565 <= lineBuffer_1564;
    end
    if (sel) begin
      lineBuffer_1566 <= lineBuffer_1565;
    end
    if (sel) begin
      lineBuffer_1567 <= lineBuffer_1566;
    end
    if (sel) begin
      lineBuffer_1568 <= lineBuffer_1567;
    end
    if (sel) begin
      lineBuffer_1569 <= lineBuffer_1568;
    end
    if (sel) begin
      lineBuffer_1570 <= lineBuffer_1569;
    end
    if (sel) begin
      lineBuffer_1571 <= lineBuffer_1570;
    end
    if (sel) begin
      lineBuffer_1572 <= lineBuffer_1571;
    end
    if (sel) begin
      lineBuffer_1573 <= lineBuffer_1572;
    end
    if (sel) begin
      lineBuffer_1574 <= lineBuffer_1573;
    end
    if (sel) begin
      lineBuffer_1575 <= lineBuffer_1574;
    end
    if (sel) begin
      lineBuffer_1576 <= lineBuffer_1575;
    end
    if (sel) begin
      lineBuffer_1577 <= lineBuffer_1576;
    end
    if (sel) begin
      lineBuffer_1578 <= lineBuffer_1577;
    end
    if (sel) begin
      lineBuffer_1579 <= lineBuffer_1578;
    end
    if (sel) begin
      lineBuffer_1580 <= lineBuffer_1579;
    end
    if (sel) begin
      lineBuffer_1581 <= lineBuffer_1580;
    end
    if (sel) begin
      lineBuffer_1582 <= lineBuffer_1581;
    end
    if (sel) begin
      lineBuffer_1583 <= lineBuffer_1582;
    end
    if (sel) begin
      lineBuffer_1584 <= lineBuffer_1583;
    end
    if (sel) begin
      lineBuffer_1585 <= lineBuffer_1584;
    end
    if (sel) begin
      lineBuffer_1586 <= lineBuffer_1585;
    end
    if (sel) begin
      lineBuffer_1587 <= lineBuffer_1586;
    end
    if (sel) begin
      lineBuffer_1588 <= lineBuffer_1587;
    end
    if (sel) begin
      lineBuffer_1589 <= lineBuffer_1588;
    end
    if (sel) begin
      lineBuffer_1590 <= lineBuffer_1589;
    end
    if (sel) begin
      lineBuffer_1591 <= lineBuffer_1590;
    end
    if (sel) begin
      lineBuffer_1592 <= lineBuffer_1591;
    end
    if (sel) begin
      lineBuffer_1593 <= lineBuffer_1592;
    end
    if (sel) begin
      lineBuffer_1594 <= lineBuffer_1593;
    end
    if (sel) begin
      lineBuffer_1595 <= lineBuffer_1594;
    end
    if (sel) begin
      lineBuffer_1596 <= lineBuffer_1595;
    end
    if (sel) begin
      lineBuffer_1597 <= lineBuffer_1596;
    end
    if (sel) begin
      lineBuffer_1598 <= lineBuffer_1597;
    end
    if (sel) begin
      lineBuffer_1599 <= lineBuffer_1598;
    end
    if (sel) begin
      lineBuffer_1600 <= lineBuffer_1599;
    end
    if (sel) begin
      lineBuffer_1601 <= lineBuffer_1600;
    end
    if (sel) begin
      lineBuffer_1602 <= lineBuffer_1601;
    end
    if (sel) begin
      lineBuffer_1603 <= lineBuffer_1602;
    end
    if (sel) begin
      lineBuffer_1604 <= lineBuffer_1603;
    end
    if (sel) begin
      lineBuffer_1605 <= lineBuffer_1604;
    end
    if (sel) begin
      lineBuffer_1606 <= lineBuffer_1605;
    end
    if (sel) begin
      lineBuffer_1607 <= lineBuffer_1606;
    end
    if (sel) begin
      lineBuffer_1608 <= lineBuffer_1607;
    end
    if (sel) begin
      lineBuffer_1609 <= lineBuffer_1608;
    end
    if (sel) begin
      lineBuffer_1610 <= lineBuffer_1609;
    end
    if (sel) begin
      lineBuffer_1611 <= lineBuffer_1610;
    end
    if (sel) begin
      lineBuffer_1612 <= lineBuffer_1611;
    end
    if (sel) begin
      lineBuffer_1613 <= lineBuffer_1612;
    end
    if (sel) begin
      lineBuffer_1614 <= lineBuffer_1613;
    end
    if (sel) begin
      lineBuffer_1615 <= lineBuffer_1614;
    end
    if (sel) begin
      lineBuffer_1616 <= lineBuffer_1615;
    end
    if (sel) begin
      lineBuffer_1617 <= lineBuffer_1616;
    end
    if (sel) begin
      lineBuffer_1618 <= lineBuffer_1617;
    end
    if (sel) begin
      lineBuffer_1619 <= lineBuffer_1618;
    end
    if (sel) begin
      lineBuffer_1620 <= lineBuffer_1619;
    end
    if (sel) begin
      lineBuffer_1621 <= lineBuffer_1620;
    end
    if (sel) begin
      lineBuffer_1622 <= lineBuffer_1621;
    end
    if (sel) begin
      lineBuffer_1623 <= lineBuffer_1622;
    end
    if (sel) begin
      lineBuffer_1624 <= lineBuffer_1623;
    end
    if (sel) begin
      lineBuffer_1625 <= lineBuffer_1624;
    end
    if (sel) begin
      lineBuffer_1626 <= lineBuffer_1625;
    end
    if (sel) begin
      lineBuffer_1627 <= lineBuffer_1626;
    end
    if (sel) begin
      lineBuffer_1628 <= lineBuffer_1627;
    end
    if (sel) begin
      lineBuffer_1629 <= lineBuffer_1628;
    end
    if (sel) begin
      lineBuffer_1630 <= lineBuffer_1629;
    end
    if (sel) begin
      lineBuffer_1631 <= lineBuffer_1630;
    end
    if (sel) begin
      lineBuffer_1632 <= lineBuffer_1631;
    end
    if (sel) begin
      lineBuffer_1633 <= lineBuffer_1632;
    end
    if (sel) begin
      lineBuffer_1634 <= lineBuffer_1633;
    end
    if (sel) begin
      lineBuffer_1635 <= lineBuffer_1634;
    end
    if (sel) begin
      lineBuffer_1636 <= lineBuffer_1635;
    end
    if (sel) begin
      lineBuffer_1637 <= lineBuffer_1636;
    end
    if (sel) begin
      lineBuffer_1638 <= lineBuffer_1637;
    end
    if (sel) begin
      lineBuffer_1639 <= lineBuffer_1638;
    end
    if (sel) begin
      lineBuffer_1640 <= lineBuffer_1639;
    end
    if (sel) begin
      lineBuffer_1641 <= lineBuffer_1640;
    end
    if (sel) begin
      lineBuffer_1642 <= lineBuffer_1641;
    end
    if (sel) begin
      lineBuffer_1643 <= lineBuffer_1642;
    end
    if (sel) begin
      lineBuffer_1644 <= lineBuffer_1643;
    end
    if (sel) begin
      lineBuffer_1645 <= lineBuffer_1644;
    end
    if (sel) begin
      lineBuffer_1646 <= lineBuffer_1645;
    end
    if (sel) begin
      lineBuffer_1647 <= lineBuffer_1646;
    end
    if (sel) begin
      lineBuffer_1648 <= lineBuffer_1647;
    end
    if (sel) begin
      lineBuffer_1649 <= lineBuffer_1648;
    end
    if (sel) begin
      lineBuffer_1650 <= lineBuffer_1649;
    end
    if (sel) begin
      lineBuffer_1651 <= lineBuffer_1650;
    end
    if (sel) begin
      lineBuffer_1652 <= lineBuffer_1651;
    end
    if (sel) begin
      lineBuffer_1653 <= lineBuffer_1652;
    end
    if (sel) begin
      lineBuffer_1654 <= lineBuffer_1653;
    end
    if (sel) begin
      lineBuffer_1655 <= lineBuffer_1654;
    end
    if (sel) begin
      lineBuffer_1656 <= lineBuffer_1655;
    end
    if (sel) begin
      lineBuffer_1657 <= lineBuffer_1656;
    end
    if (sel) begin
      lineBuffer_1658 <= lineBuffer_1657;
    end
    if (sel) begin
      lineBuffer_1659 <= lineBuffer_1658;
    end
    if (sel) begin
      lineBuffer_1660 <= lineBuffer_1659;
    end
    if (sel) begin
      lineBuffer_1661 <= lineBuffer_1660;
    end
    if (sel) begin
      lineBuffer_1662 <= lineBuffer_1661;
    end
    if (sel) begin
      lineBuffer_1663 <= lineBuffer_1662;
    end
    if (sel) begin
      lineBuffer_1664 <= lineBuffer_1663;
    end
    if (sel) begin
      lineBuffer_1665 <= lineBuffer_1664;
    end
    if (sel) begin
      lineBuffer_1666 <= lineBuffer_1665;
    end
    if (sel) begin
      lineBuffer_1667 <= lineBuffer_1666;
    end
    if (sel) begin
      lineBuffer_1668 <= lineBuffer_1667;
    end
    if (sel) begin
      lineBuffer_1669 <= lineBuffer_1668;
    end
    if (sel) begin
      lineBuffer_1670 <= lineBuffer_1669;
    end
    if (sel) begin
      lineBuffer_1671 <= lineBuffer_1670;
    end
    if (sel) begin
      lineBuffer_1672 <= lineBuffer_1671;
    end
    if (sel) begin
      lineBuffer_1673 <= lineBuffer_1672;
    end
    if (sel) begin
      lineBuffer_1674 <= lineBuffer_1673;
    end
    if (sel) begin
      lineBuffer_1675 <= lineBuffer_1674;
    end
    if (sel) begin
      lineBuffer_1676 <= lineBuffer_1675;
    end
    if (sel) begin
      lineBuffer_1677 <= lineBuffer_1676;
    end
    if (sel) begin
      lineBuffer_1678 <= lineBuffer_1677;
    end
    if (sel) begin
      lineBuffer_1679 <= lineBuffer_1678;
    end
    if (sel) begin
      lineBuffer_1680 <= lineBuffer_1679;
    end
    if (sel) begin
      lineBuffer_1681 <= lineBuffer_1680;
    end
    if (sel) begin
      lineBuffer_1682 <= lineBuffer_1681;
    end
    if (sel) begin
      lineBuffer_1683 <= lineBuffer_1682;
    end
    if (sel) begin
      lineBuffer_1684 <= lineBuffer_1683;
    end
    if (sel) begin
      lineBuffer_1685 <= lineBuffer_1684;
    end
    if (sel) begin
      lineBuffer_1686 <= lineBuffer_1685;
    end
    if (sel) begin
      lineBuffer_1687 <= lineBuffer_1686;
    end
    if (sel) begin
      lineBuffer_1688 <= lineBuffer_1687;
    end
    if (sel) begin
      lineBuffer_1689 <= lineBuffer_1688;
    end
    if (sel) begin
      lineBuffer_1690 <= lineBuffer_1689;
    end
    if (sel) begin
      lineBuffer_1691 <= lineBuffer_1690;
    end
    if (sel) begin
      lineBuffer_1692 <= lineBuffer_1691;
    end
    if (sel) begin
      lineBuffer_1693 <= lineBuffer_1692;
    end
    if (sel) begin
      lineBuffer_1694 <= lineBuffer_1693;
    end
    if (sel) begin
      lineBuffer_1695 <= lineBuffer_1694;
    end
    if (sel) begin
      lineBuffer_1696 <= lineBuffer_1695;
    end
    if (sel) begin
      lineBuffer_1697 <= lineBuffer_1696;
    end
    if (sel) begin
      lineBuffer_1698 <= lineBuffer_1697;
    end
    if (sel) begin
      lineBuffer_1699 <= lineBuffer_1698;
    end
    if (sel) begin
      lineBuffer_1700 <= lineBuffer_1699;
    end
    if (sel) begin
      lineBuffer_1701 <= lineBuffer_1700;
    end
    if (sel) begin
      lineBuffer_1702 <= lineBuffer_1701;
    end
    if (sel) begin
      lineBuffer_1703 <= lineBuffer_1702;
    end
    if (sel) begin
      lineBuffer_1704 <= lineBuffer_1703;
    end
    if (sel) begin
      lineBuffer_1705 <= lineBuffer_1704;
    end
    if (sel) begin
      lineBuffer_1706 <= lineBuffer_1705;
    end
    if (sel) begin
      lineBuffer_1707 <= lineBuffer_1706;
    end
    if (sel) begin
      lineBuffer_1708 <= lineBuffer_1707;
    end
    if (sel) begin
      lineBuffer_1709 <= lineBuffer_1708;
    end
    if (sel) begin
      lineBuffer_1710 <= lineBuffer_1709;
    end
    if (sel) begin
      lineBuffer_1711 <= lineBuffer_1710;
    end
    if (sel) begin
      lineBuffer_1712 <= lineBuffer_1711;
    end
    if (sel) begin
      lineBuffer_1713 <= lineBuffer_1712;
    end
    if (sel) begin
      lineBuffer_1714 <= lineBuffer_1713;
    end
    if (sel) begin
      lineBuffer_1715 <= lineBuffer_1714;
    end
    if (sel) begin
      lineBuffer_1716 <= lineBuffer_1715;
    end
    if (sel) begin
      lineBuffer_1717 <= lineBuffer_1716;
    end
    if (sel) begin
      lineBuffer_1718 <= lineBuffer_1717;
    end
    if (sel) begin
      lineBuffer_1719 <= lineBuffer_1718;
    end
    if (sel) begin
      lineBuffer_1720 <= lineBuffer_1719;
    end
    if (sel) begin
      lineBuffer_1721 <= lineBuffer_1720;
    end
    if (sel) begin
      lineBuffer_1722 <= lineBuffer_1721;
    end
    if (sel) begin
      lineBuffer_1723 <= lineBuffer_1722;
    end
    if (sel) begin
      lineBuffer_1724 <= lineBuffer_1723;
    end
    if (sel) begin
      lineBuffer_1725 <= lineBuffer_1724;
    end
    if (sel) begin
      lineBuffer_1726 <= lineBuffer_1725;
    end
    if (sel) begin
      lineBuffer_1727 <= lineBuffer_1726;
    end
    if (sel) begin
      lineBuffer_1728 <= lineBuffer_1727;
    end
    if (sel) begin
      lineBuffer_1729 <= lineBuffer_1728;
    end
    if (sel) begin
      lineBuffer_1730 <= lineBuffer_1729;
    end
    if (sel) begin
      lineBuffer_1731 <= lineBuffer_1730;
    end
    if (sel) begin
      lineBuffer_1732 <= lineBuffer_1731;
    end
    if (sel) begin
      lineBuffer_1733 <= lineBuffer_1732;
    end
    if (sel) begin
      lineBuffer_1734 <= lineBuffer_1733;
    end
    if (sel) begin
      lineBuffer_1735 <= lineBuffer_1734;
    end
    if (sel) begin
      lineBuffer_1736 <= lineBuffer_1735;
    end
    if (sel) begin
      lineBuffer_1737 <= lineBuffer_1736;
    end
    if (sel) begin
      lineBuffer_1738 <= lineBuffer_1737;
    end
    if (sel) begin
      lineBuffer_1739 <= lineBuffer_1738;
    end
    if (sel) begin
      lineBuffer_1740 <= lineBuffer_1739;
    end
    if (sel) begin
      lineBuffer_1741 <= lineBuffer_1740;
    end
    if (sel) begin
      lineBuffer_1742 <= lineBuffer_1741;
    end
    if (sel) begin
      lineBuffer_1743 <= lineBuffer_1742;
    end
    if (sel) begin
      lineBuffer_1744 <= lineBuffer_1743;
    end
    if (sel) begin
      lineBuffer_1745 <= lineBuffer_1744;
    end
    if (sel) begin
      lineBuffer_1746 <= lineBuffer_1745;
    end
    if (sel) begin
      lineBuffer_1747 <= lineBuffer_1746;
    end
    if (sel) begin
      lineBuffer_1748 <= lineBuffer_1747;
    end
    if (sel) begin
      lineBuffer_1749 <= lineBuffer_1748;
    end
    if (sel) begin
      lineBuffer_1750 <= lineBuffer_1749;
    end
    if (sel) begin
      lineBuffer_1751 <= lineBuffer_1750;
    end
    if (sel) begin
      lineBuffer_1752 <= lineBuffer_1751;
    end
    if (sel) begin
      lineBuffer_1753 <= lineBuffer_1752;
    end
    if (sel) begin
      lineBuffer_1754 <= lineBuffer_1753;
    end
    if (sel) begin
      lineBuffer_1755 <= lineBuffer_1754;
    end
    if (sel) begin
      lineBuffer_1756 <= lineBuffer_1755;
    end
    if (sel) begin
      lineBuffer_1757 <= lineBuffer_1756;
    end
    if (sel) begin
      lineBuffer_1758 <= lineBuffer_1757;
    end
    if (sel) begin
      lineBuffer_1759 <= lineBuffer_1758;
    end
    if (sel) begin
      lineBuffer_1760 <= lineBuffer_1759;
    end
    if (sel) begin
      lineBuffer_1761 <= lineBuffer_1760;
    end
    if (sel) begin
      lineBuffer_1762 <= lineBuffer_1761;
    end
    if (sel) begin
      lineBuffer_1763 <= lineBuffer_1762;
    end
    if (sel) begin
      lineBuffer_1764 <= lineBuffer_1763;
    end
    if (sel) begin
      lineBuffer_1765 <= lineBuffer_1764;
    end
    if (sel) begin
      lineBuffer_1766 <= lineBuffer_1765;
    end
    if (sel) begin
      lineBuffer_1767 <= lineBuffer_1766;
    end
    if (sel) begin
      lineBuffer_1768 <= lineBuffer_1767;
    end
    if (sel) begin
      lineBuffer_1769 <= lineBuffer_1768;
    end
    if (sel) begin
      lineBuffer_1770 <= lineBuffer_1769;
    end
    if (sel) begin
      lineBuffer_1771 <= lineBuffer_1770;
    end
    if (sel) begin
      lineBuffer_1772 <= lineBuffer_1771;
    end
    if (sel) begin
      lineBuffer_1773 <= lineBuffer_1772;
    end
    if (sel) begin
      lineBuffer_1774 <= lineBuffer_1773;
    end
    if (sel) begin
      lineBuffer_1775 <= lineBuffer_1774;
    end
    if (sel) begin
      lineBuffer_1776 <= lineBuffer_1775;
    end
    if (sel) begin
      lineBuffer_1777 <= lineBuffer_1776;
    end
    if (sel) begin
      lineBuffer_1778 <= lineBuffer_1777;
    end
    if (sel) begin
      lineBuffer_1779 <= lineBuffer_1778;
    end
    if (sel) begin
      lineBuffer_1780 <= lineBuffer_1779;
    end
    if (sel) begin
      lineBuffer_1781 <= lineBuffer_1780;
    end
    if (sel) begin
      lineBuffer_1782 <= lineBuffer_1781;
    end
    if (sel) begin
      lineBuffer_1783 <= lineBuffer_1782;
    end
    if (sel) begin
      lineBuffer_1784 <= lineBuffer_1783;
    end
    if (sel) begin
      lineBuffer_1785 <= lineBuffer_1784;
    end
    if (sel) begin
      lineBuffer_1786 <= lineBuffer_1785;
    end
    if (sel) begin
      lineBuffer_1787 <= lineBuffer_1786;
    end
    if (sel) begin
      lineBuffer_1788 <= lineBuffer_1787;
    end
    if (sel) begin
      lineBuffer_1789 <= lineBuffer_1788;
    end
    if (sel) begin
      lineBuffer_1790 <= lineBuffer_1789;
    end
    if (sel) begin
      lineBuffer_1791 <= lineBuffer_1790;
    end
    if (sel) begin
      lineBuffer_1792 <= lineBuffer_1791;
    end
    if (sel) begin
      lineBuffer_1793 <= lineBuffer_1792;
    end
    if (sel) begin
      lineBuffer_1794 <= lineBuffer_1793;
    end
    if (sel) begin
      lineBuffer_1795 <= lineBuffer_1794;
    end
    if (sel) begin
      lineBuffer_1796 <= lineBuffer_1795;
    end
    if (sel) begin
      lineBuffer_1797 <= lineBuffer_1796;
    end
    if (sel) begin
      lineBuffer_1798 <= lineBuffer_1797;
    end
    if (sel) begin
      lineBuffer_1799 <= lineBuffer_1798;
    end
    if (sel) begin
      lineBuffer_1800 <= lineBuffer_1799;
    end
    if (sel) begin
      lineBuffer_1801 <= lineBuffer_1800;
    end
    if (sel) begin
      lineBuffer_1802 <= lineBuffer_1801;
    end
    if (sel) begin
      lineBuffer_1803 <= lineBuffer_1802;
    end
    if (sel) begin
      lineBuffer_1804 <= lineBuffer_1803;
    end
    if (sel) begin
      lineBuffer_1805 <= lineBuffer_1804;
    end
    if (sel) begin
      lineBuffer_1806 <= lineBuffer_1805;
    end
    if (sel) begin
      lineBuffer_1807 <= lineBuffer_1806;
    end
    if (sel) begin
      lineBuffer_1808 <= lineBuffer_1807;
    end
    if (sel) begin
      lineBuffer_1809 <= lineBuffer_1808;
    end
    if (sel) begin
      lineBuffer_1810 <= lineBuffer_1809;
    end
    if (sel) begin
      lineBuffer_1811 <= lineBuffer_1810;
    end
    if (sel) begin
      lineBuffer_1812 <= lineBuffer_1811;
    end
    if (sel) begin
      lineBuffer_1813 <= lineBuffer_1812;
    end
    if (sel) begin
      lineBuffer_1814 <= lineBuffer_1813;
    end
    if (sel) begin
      lineBuffer_1815 <= lineBuffer_1814;
    end
    if (sel) begin
      lineBuffer_1816 <= lineBuffer_1815;
    end
    if (sel) begin
      lineBuffer_1817 <= lineBuffer_1816;
    end
    if (sel) begin
      lineBuffer_1818 <= lineBuffer_1817;
    end
    if (sel) begin
      lineBuffer_1819 <= lineBuffer_1818;
    end
    if (sel) begin
      lineBuffer_1820 <= lineBuffer_1819;
    end
    if (sel) begin
      lineBuffer_1821 <= lineBuffer_1820;
    end
    if (sel) begin
      lineBuffer_1822 <= lineBuffer_1821;
    end
    if (sel) begin
      lineBuffer_1823 <= lineBuffer_1822;
    end
    if (sel) begin
      lineBuffer_1824 <= lineBuffer_1823;
    end
    if (sel) begin
      lineBuffer_1825 <= lineBuffer_1824;
    end
    if (sel) begin
      lineBuffer_1826 <= lineBuffer_1825;
    end
    if (sel) begin
      lineBuffer_1827 <= lineBuffer_1826;
    end
    if (sel) begin
      lineBuffer_1828 <= lineBuffer_1827;
    end
    if (sel) begin
      lineBuffer_1829 <= lineBuffer_1828;
    end
    if (sel) begin
      lineBuffer_1830 <= lineBuffer_1829;
    end
    if (sel) begin
      lineBuffer_1831 <= lineBuffer_1830;
    end
    if (sel) begin
      lineBuffer_1832 <= lineBuffer_1831;
    end
    if (sel) begin
      lineBuffer_1833 <= lineBuffer_1832;
    end
    if (sel) begin
      lineBuffer_1834 <= lineBuffer_1833;
    end
    if (sel) begin
      lineBuffer_1835 <= lineBuffer_1834;
    end
    if (sel) begin
      lineBuffer_1836 <= lineBuffer_1835;
    end
    if (sel) begin
      lineBuffer_1837 <= lineBuffer_1836;
    end
    if (sel) begin
      lineBuffer_1838 <= lineBuffer_1837;
    end
    if (sel) begin
      lineBuffer_1839 <= lineBuffer_1838;
    end
    if (sel) begin
      lineBuffer_1840 <= lineBuffer_1839;
    end
    if (sel) begin
      lineBuffer_1841 <= lineBuffer_1840;
    end
    if (sel) begin
      lineBuffer_1842 <= lineBuffer_1841;
    end
    if (sel) begin
      lineBuffer_1843 <= lineBuffer_1842;
    end
    if (sel) begin
      lineBuffer_1844 <= lineBuffer_1843;
    end
    if (sel) begin
      lineBuffer_1845 <= lineBuffer_1844;
    end
    if (sel) begin
      lineBuffer_1846 <= lineBuffer_1845;
    end
    if (sel) begin
      lineBuffer_1847 <= lineBuffer_1846;
    end
    if (sel) begin
      lineBuffer_1848 <= lineBuffer_1847;
    end
    if (sel) begin
      lineBuffer_1849 <= lineBuffer_1848;
    end
    if (sel) begin
      lineBuffer_1850 <= lineBuffer_1849;
    end
    if (sel) begin
      lineBuffer_1851 <= lineBuffer_1850;
    end
    if (sel) begin
      lineBuffer_1852 <= lineBuffer_1851;
    end
    if (sel) begin
      lineBuffer_1853 <= lineBuffer_1852;
    end
    if (sel) begin
      lineBuffer_1854 <= lineBuffer_1853;
    end
    if (sel) begin
      lineBuffer_1855 <= lineBuffer_1854;
    end
    if (sel) begin
      lineBuffer_1856 <= lineBuffer_1855;
    end
    if (sel) begin
      lineBuffer_1857 <= lineBuffer_1856;
    end
    if (sel) begin
      lineBuffer_1858 <= lineBuffer_1857;
    end
    if (sel) begin
      lineBuffer_1859 <= lineBuffer_1858;
    end
    if (sel) begin
      lineBuffer_1860 <= lineBuffer_1859;
    end
    if (sel) begin
      lineBuffer_1861 <= lineBuffer_1860;
    end
    if (sel) begin
      lineBuffer_1862 <= lineBuffer_1861;
    end
    if (sel) begin
      lineBuffer_1863 <= lineBuffer_1862;
    end
    if (sel) begin
      lineBuffer_1864 <= lineBuffer_1863;
    end
    if (sel) begin
      lineBuffer_1865 <= lineBuffer_1864;
    end
    if (sel) begin
      lineBuffer_1866 <= lineBuffer_1865;
    end
    if (sel) begin
      lineBuffer_1867 <= lineBuffer_1866;
    end
    if (sel) begin
      lineBuffer_1868 <= lineBuffer_1867;
    end
    if (sel) begin
      lineBuffer_1869 <= lineBuffer_1868;
    end
    if (sel) begin
      lineBuffer_1870 <= lineBuffer_1869;
    end
    if (sel) begin
      lineBuffer_1871 <= lineBuffer_1870;
    end
    if (sel) begin
      lineBuffer_1872 <= lineBuffer_1871;
    end
    if (sel) begin
      lineBuffer_1873 <= lineBuffer_1872;
    end
    if (sel) begin
      lineBuffer_1874 <= lineBuffer_1873;
    end
    if (sel) begin
      lineBuffer_1875 <= lineBuffer_1874;
    end
    if (sel) begin
      lineBuffer_1876 <= lineBuffer_1875;
    end
    if (sel) begin
      lineBuffer_1877 <= lineBuffer_1876;
    end
    if (sel) begin
      lineBuffer_1878 <= lineBuffer_1877;
    end
    if (sel) begin
      lineBuffer_1879 <= lineBuffer_1878;
    end
    if (sel) begin
      lineBuffer_1880 <= lineBuffer_1879;
    end
    if (sel) begin
      lineBuffer_1881 <= lineBuffer_1880;
    end
    if (sel) begin
      lineBuffer_1882 <= lineBuffer_1881;
    end
    if (sel) begin
      lineBuffer_1883 <= lineBuffer_1882;
    end
    if (sel) begin
      lineBuffer_1884 <= lineBuffer_1883;
    end
    if (sel) begin
      lineBuffer_1885 <= lineBuffer_1884;
    end
    if (sel) begin
      lineBuffer_1886 <= lineBuffer_1885;
    end
    if (sel) begin
      lineBuffer_1887 <= lineBuffer_1886;
    end
    if (sel) begin
      lineBuffer_1888 <= lineBuffer_1887;
    end
    if (sel) begin
      lineBuffer_1889 <= lineBuffer_1888;
    end
    if (sel) begin
      lineBuffer_1890 <= lineBuffer_1889;
    end
    if (sel) begin
      lineBuffer_1891 <= lineBuffer_1890;
    end
    if (sel) begin
      lineBuffer_1892 <= lineBuffer_1891;
    end
    if (sel) begin
      lineBuffer_1893 <= lineBuffer_1892;
    end
    if (sel) begin
      lineBuffer_1894 <= lineBuffer_1893;
    end
    if (sel) begin
      lineBuffer_1895 <= lineBuffer_1894;
    end
    if (sel) begin
      lineBuffer_1896 <= lineBuffer_1895;
    end
    if (sel) begin
      lineBuffer_1897 <= lineBuffer_1896;
    end
    if (sel) begin
      lineBuffer_1898 <= lineBuffer_1897;
    end
    if (sel) begin
      lineBuffer_1899 <= lineBuffer_1898;
    end
    if (sel) begin
      lineBuffer_1900 <= lineBuffer_1899;
    end
    if (sel) begin
      lineBuffer_1901 <= lineBuffer_1900;
    end
    if (sel) begin
      lineBuffer_1902 <= lineBuffer_1901;
    end
    if (sel) begin
      lineBuffer_1903 <= lineBuffer_1902;
    end
    if (sel) begin
      lineBuffer_1904 <= lineBuffer_1903;
    end
    if (sel) begin
      lineBuffer_1905 <= lineBuffer_1904;
    end
    if (sel) begin
      lineBuffer_1906 <= lineBuffer_1905;
    end
    if (sel) begin
      lineBuffer_1907 <= lineBuffer_1906;
    end
    if (sel) begin
      lineBuffer_1908 <= lineBuffer_1907;
    end
    if (sel) begin
      lineBuffer_1909 <= lineBuffer_1908;
    end
    if (sel) begin
      lineBuffer_1910 <= lineBuffer_1909;
    end
    if (sel) begin
      lineBuffer_1911 <= lineBuffer_1910;
    end
    if (sel) begin
      lineBuffer_1912 <= lineBuffer_1911;
    end
    if (sel) begin
      lineBuffer_1913 <= lineBuffer_1912;
    end
    if (sel) begin
      lineBuffer_1914 <= lineBuffer_1913;
    end
    if (sel) begin
      lineBuffer_1915 <= lineBuffer_1914;
    end
    if (sel) begin
      lineBuffer_1916 <= lineBuffer_1915;
    end
    if (sel) begin
      lineBuffer_1917 <= lineBuffer_1916;
    end
    if (sel) begin
      lineBuffer_1918 <= lineBuffer_1917;
    end
    if (sel) begin
      lineBuffer_1919 <= lineBuffer_1918;
    end
    if (sel) begin
      lineBuffer_1920 <= lineBuffer_1919;
    end
    if (sel) begin
      lineBuffer_1921 <= lineBuffer_1920;
    end
    if (sel) begin
      lineBuffer_1922 <= lineBuffer_1921;
    end
    if (sel) begin
      lineBuffer_1923 <= lineBuffer_1922;
    end
    if (sel) begin
      lineBuffer_1924 <= lineBuffer_1923;
    end
    if (sel) begin
      lineBuffer_1925 <= lineBuffer_1924;
    end
    if (sel) begin
      lineBuffer_1926 <= lineBuffer_1925;
    end
    if (sel) begin
      lineBuffer_1927 <= lineBuffer_1926;
    end
    if (sel) begin
      lineBuffer_1928 <= lineBuffer_1927;
    end
    if (sel) begin
      lineBuffer_1929 <= lineBuffer_1928;
    end
    if (sel) begin
      lineBuffer_1930 <= lineBuffer_1929;
    end
    if (sel) begin
      lineBuffer_1931 <= lineBuffer_1930;
    end
    if (sel) begin
      lineBuffer_1932 <= lineBuffer_1931;
    end
    if (sel) begin
      lineBuffer_1933 <= lineBuffer_1932;
    end
    if (sel) begin
      lineBuffer_1934 <= lineBuffer_1933;
    end
    if (sel) begin
      lineBuffer_1935 <= lineBuffer_1934;
    end
    if (sel) begin
      lineBuffer_1936 <= lineBuffer_1935;
    end
    if (sel) begin
      lineBuffer_1937 <= lineBuffer_1936;
    end
    if (sel) begin
      lineBuffer_1938 <= lineBuffer_1937;
    end
    if (sel) begin
      lineBuffer_1939 <= lineBuffer_1938;
    end
    if (sel) begin
      lineBuffer_1940 <= lineBuffer_1939;
    end
    if (sel) begin
      lineBuffer_1941 <= lineBuffer_1940;
    end
    if (sel) begin
      lineBuffer_1942 <= lineBuffer_1941;
    end
    if (sel) begin
      lineBuffer_1943 <= lineBuffer_1942;
    end
    if (sel) begin
      lineBuffer_1944 <= lineBuffer_1943;
    end
    if (sel) begin
      lineBuffer_1945 <= lineBuffer_1944;
    end
    if (sel) begin
      lineBuffer_1946 <= lineBuffer_1945;
    end
    if (sel) begin
      lineBuffer_1947 <= lineBuffer_1946;
    end
    if (sel) begin
      lineBuffer_1948 <= lineBuffer_1947;
    end
    if (sel) begin
      lineBuffer_1949 <= lineBuffer_1948;
    end
    if (sel) begin
      lineBuffer_1950 <= lineBuffer_1949;
    end
    if (sel) begin
      lineBuffer_1951 <= lineBuffer_1950;
    end
    if (sel) begin
      lineBuffer_1952 <= lineBuffer_1951;
    end
    if (sel) begin
      lineBuffer_1953 <= lineBuffer_1952;
    end
    if (sel) begin
      lineBuffer_1954 <= lineBuffer_1953;
    end
    if (sel) begin
      lineBuffer_1955 <= lineBuffer_1954;
    end
    if (sel) begin
      lineBuffer_1956 <= lineBuffer_1955;
    end
    if (sel) begin
      lineBuffer_1957 <= lineBuffer_1956;
    end
    if (sel) begin
      lineBuffer_1958 <= lineBuffer_1957;
    end
    if (sel) begin
      lineBuffer_1959 <= lineBuffer_1958;
    end
    if (sel) begin
      lineBuffer_1960 <= lineBuffer_1959;
    end
    if (sel) begin
      lineBuffer_1961 <= lineBuffer_1960;
    end
    if (sel) begin
      lineBuffer_1962 <= lineBuffer_1961;
    end
    if (sel) begin
      lineBuffer_1963 <= lineBuffer_1962;
    end
    if (sel) begin
      lineBuffer_1964 <= lineBuffer_1963;
    end
    if (sel) begin
      lineBuffer_1965 <= lineBuffer_1964;
    end
    if (sel) begin
      lineBuffer_1966 <= lineBuffer_1965;
    end
    if (sel) begin
      lineBuffer_1967 <= lineBuffer_1966;
    end
    if (sel) begin
      lineBuffer_1968 <= lineBuffer_1967;
    end
    if (sel) begin
      lineBuffer_1969 <= lineBuffer_1968;
    end
    if (sel) begin
      lineBuffer_1970 <= lineBuffer_1969;
    end
    if (sel) begin
      lineBuffer_1971 <= lineBuffer_1970;
    end
    if (sel) begin
      lineBuffer_1972 <= lineBuffer_1971;
    end
    if (sel) begin
      lineBuffer_1973 <= lineBuffer_1972;
    end
    if (sel) begin
      lineBuffer_1974 <= lineBuffer_1973;
    end
    if (sel) begin
      lineBuffer_1975 <= lineBuffer_1974;
    end
    if (sel) begin
      lineBuffer_1976 <= lineBuffer_1975;
    end
    if (sel) begin
      lineBuffer_1977 <= lineBuffer_1976;
    end
    if (sel) begin
      lineBuffer_1978 <= lineBuffer_1977;
    end
    if (sel) begin
      lineBuffer_1979 <= lineBuffer_1978;
    end
    if (sel) begin
      lineBuffer_1980 <= lineBuffer_1979;
    end
    if (sel) begin
      lineBuffer_1981 <= lineBuffer_1980;
    end
    if (sel) begin
      lineBuffer_1982 <= lineBuffer_1981;
    end
    if (sel) begin
      lineBuffer_1983 <= lineBuffer_1982;
    end
    if (sel) begin
      lineBuffer_1984 <= lineBuffer_1983;
    end
    if (sel) begin
      lineBuffer_1985 <= lineBuffer_1984;
    end
    if (sel) begin
      lineBuffer_1986 <= lineBuffer_1985;
    end
    if (sel) begin
      lineBuffer_1987 <= lineBuffer_1986;
    end
    if (sel) begin
      lineBuffer_1988 <= lineBuffer_1987;
    end
    if (sel) begin
      lineBuffer_1989 <= lineBuffer_1988;
    end
    if (sel) begin
      lineBuffer_1990 <= lineBuffer_1989;
    end
    if (sel) begin
      lineBuffer_1991 <= lineBuffer_1990;
    end
    if (sel) begin
      lineBuffer_1992 <= lineBuffer_1991;
    end
    if (sel) begin
      lineBuffer_1993 <= lineBuffer_1992;
    end
    if (sel) begin
      lineBuffer_1994 <= lineBuffer_1993;
    end
    if (sel) begin
      lineBuffer_1995 <= lineBuffer_1994;
    end
    if (sel) begin
      lineBuffer_1996 <= lineBuffer_1995;
    end
    if (sel) begin
      lineBuffer_1997 <= lineBuffer_1996;
    end
    if (sel) begin
      lineBuffer_1998 <= lineBuffer_1997;
    end
    if (sel) begin
      lineBuffer_1999 <= lineBuffer_1998;
    end
    if (sel) begin
      lineBuffer_2000 <= lineBuffer_1999;
    end
    if (sel) begin
      lineBuffer_2001 <= lineBuffer_2000;
    end
    if (sel) begin
      lineBuffer_2002 <= lineBuffer_2001;
    end
    if (sel) begin
      lineBuffer_2003 <= lineBuffer_2002;
    end
    if (sel) begin
      lineBuffer_2004 <= lineBuffer_2003;
    end
    if (sel) begin
      lineBuffer_2005 <= lineBuffer_2004;
    end
    if (sel) begin
      lineBuffer_2006 <= lineBuffer_2005;
    end
    if (sel) begin
      lineBuffer_2007 <= lineBuffer_2006;
    end
    if (sel) begin
      lineBuffer_2008 <= lineBuffer_2007;
    end
    if (sel) begin
      lineBuffer_2009 <= lineBuffer_2008;
    end
    if (sel) begin
      lineBuffer_2010 <= lineBuffer_2009;
    end
    if (sel) begin
      lineBuffer_2011 <= lineBuffer_2010;
    end
    if (sel) begin
      lineBuffer_2012 <= lineBuffer_2011;
    end
    if (sel) begin
      lineBuffer_2013 <= lineBuffer_2012;
    end
    if (sel) begin
      lineBuffer_2014 <= lineBuffer_2013;
    end
    if (sel) begin
      lineBuffer_2015 <= lineBuffer_2014;
    end
    if (sel) begin
      lineBuffer_2016 <= lineBuffer_2015;
    end
    if (sel) begin
      lineBuffer_2017 <= lineBuffer_2016;
    end
    if (sel) begin
      lineBuffer_2018 <= lineBuffer_2017;
    end
    if (sel) begin
      lineBuffer_2019 <= lineBuffer_2018;
    end
    if (sel) begin
      lineBuffer_2020 <= lineBuffer_2019;
    end
    if (sel) begin
      lineBuffer_2021 <= lineBuffer_2020;
    end
    if (sel) begin
      lineBuffer_2022 <= lineBuffer_2021;
    end
    if (sel) begin
      lineBuffer_2023 <= lineBuffer_2022;
    end
    if (sel) begin
      lineBuffer_2024 <= lineBuffer_2023;
    end
    if (sel) begin
      lineBuffer_2025 <= lineBuffer_2024;
    end
    if (sel) begin
      lineBuffer_2026 <= lineBuffer_2025;
    end
    if (sel) begin
      lineBuffer_2027 <= lineBuffer_2026;
    end
    if (sel) begin
      lineBuffer_2028 <= lineBuffer_2027;
    end
    if (sel) begin
      lineBuffer_2029 <= lineBuffer_2028;
    end
    if (sel) begin
      lineBuffer_2030 <= lineBuffer_2029;
    end
    if (sel) begin
      lineBuffer_2031 <= lineBuffer_2030;
    end
    if (sel) begin
      lineBuffer_2032 <= lineBuffer_2031;
    end
    if (sel) begin
      lineBuffer_2033 <= lineBuffer_2032;
    end
    if (sel) begin
      lineBuffer_2034 <= lineBuffer_2033;
    end
    if (sel) begin
      lineBuffer_2035 <= lineBuffer_2034;
    end
    if (sel) begin
      lineBuffer_2036 <= lineBuffer_2035;
    end
    if (sel) begin
      lineBuffer_2037 <= lineBuffer_2036;
    end
    if (sel) begin
      lineBuffer_2038 <= lineBuffer_2037;
    end
    if (sel) begin
      lineBuffer_2039 <= lineBuffer_2038;
    end
    if (sel) begin
      lineBuffer_2040 <= lineBuffer_2039;
    end
    if (sel) begin
      lineBuffer_2041 <= lineBuffer_2040;
    end
    if (sel) begin
      lineBuffer_2042 <= lineBuffer_2041;
    end
    if (sel) begin
      lineBuffer_2043 <= lineBuffer_2042;
    end
    if (sel) begin
      lineBuffer_2044 <= lineBuffer_2043;
    end
    if (sel) begin
      lineBuffer_2045 <= lineBuffer_2044;
    end
    if (sel) begin
      lineBuffer_2046 <= lineBuffer_2045;
    end
    if (sel) begin
      lineBuffer_2047 <= lineBuffer_2046;
    end
    if (sel) begin
      lineBuffer_2048 <= lineBuffer_2047;
    end
    if (sel) begin
      lineBuffer_2049 <= lineBuffer_2048;
    end
    if (sel) begin
      lineBuffer_2050 <= lineBuffer_2049;
    end
    if (sel) begin
      lineBuffer_2051 <= lineBuffer_2050;
    end
    if (sel) begin
      lineBuffer_2052 <= lineBuffer_2051;
    end
    if (sel) begin
      lineBuffer_2053 <= lineBuffer_2052;
    end
    if (sel) begin
      lineBuffer_2054 <= lineBuffer_2053;
    end
    if (sel) begin
      lineBuffer_2055 <= lineBuffer_2054;
    end
    if (sel) begin
      lineBuffer_2056 <= lineBuffer_2055;
    end
    if (sel) begin
      lineBuffer_2057 <= lineBuffer_2056;
    end
    if (sel) begin
      lineBuffer_2058 <= lineBuffer_2057;
    end
    if (sel) begin
      lineBuffer_2059 <= lineBuffer_2058;
    end
    if (sel) begin
      lineBuffer_2060 <= lineBuffer_2059;
    end
    if (sel) begin
      lineBuffer_2061 <= lineBuffer_2060;
    end
    if (sel) begin
      lineBuffer_2062 <= lineBuffer_2061;
    end
    if (sel) begin
      lineBuffer_2063 <= lineBuffer_2062;
    end
    if (sel) begin
      lineBuffer_2064 <= lineBuffer_2063;
    end
    if (sel) begin
      lineBuffer_2065 <= lineBuffer_2064;
    end
    if (sel) begin
      lineBuffer_2066 <= lineBuffer_2065;
    end
    if (sel) begin
      lineBuffer_2067 <= lineBuffer_2066;
    end
    if (sel) begin
      lineBuffer_2068 <= lineBuffer_2067;
    end
    if (sel) begin
      lineBuffer_2069 <= lineBuffer_2068;
    end
    if (sel) begin
      lineBuffer_2070 <= lineBuffer_2069;
    end
    if (sel) begin
      lineBuffer_2071 <= lineBuffer_2070;
    end
    if (sel) begin
      lineBuffer_2072 <= lineBuffer_2071;
    end
    if (sel) begin
      lineBuffer_2073 <= lineBuffer_2072;
    end
    if (sel) begin
      lineBuffer_2074 <= lineBuffer_2073;
    end
    if (sel) begin
      lineBuffer_2075 <= lineBuffer_2074;
    end
    if (sel) begin
      lineBuffer_2076 <= lineBuffer_2075;
    end
    if (sel) begin
      lineBuffer_2077 <= lineBuffer_2076;
    end
    if (sel) begin
      lineBuffer_2078 <= lineBuffer_2077;
    end
    if (sel) begin
      lineBuffer_2079 <= lineBuffer_2078;
    end
    if (sel) begin
      lineBuffer_2080 <= lineBuffer_2079;
    end
    if (sel) begin
      lineBuffer_2081 <= lineBuffer_2080;
    end
    if (sel) begin
      lineBuffer_2082 <= lineBuffer_2081;
    end
    if (sel) begin
      lineBuffer_2083 <= lineBuffer_2082;
    end
    if (sel) begin
      lineBuffer_2084 <= lineBuffer_2083;
    end
    if (sel) begin
      lineBuffer_2085 <= lineBuffer_2084;
    end
    if (sel) begin
      lineBuffer_2086 <= lineBuffer_2085;
    end
    if (sel) begin
      lineBuffer_2087 <= lineBuffer_2086;
    end
    if (sel) begin
      lineBuffer_2088 <= lineBuffer_2087;
    end
    if (sel) begin
      lineBuffer_2089 <= lineBuffer_2088;
    end
    if (sel) begin
      lineBuffer_2090 <= lineBuffer_2089;
    end
    if (sel) begin
      lineBuffer_2091 <= lineBuffer_2090;
    end
    if (sel) begin
      lineBuffer_2092 <= lineBuffer_2091;
    end
    if (sel) begin
      lineBuffer_2093 <= lineBuffer_2092;
    end
    if (sel) begin
      lineBuffer_2094 <= lineBuffer_2093;
    end
    if (sel) begin
      lineBuffer_2095 <= lineBuffer_2094;
    end
    if (sel) begin
      lineBuffer_2096 <= lineBuffer_2095;
    end
    if (sel) begin
      lineBuffer_2097 <= lineBuffer_2096;
    end
    if (sel) begin
      lineBuffer_2098 <= lineBuffer_2097;
    end
    if (sel) begin
      lineBuffer_2099 <= lineBuffer_2098;
    end
    if (sel) begin
      lineBuffer_2100 <= lineBuffer_2099;
    end
    if (sel) begin
      lineBuffer_2101 <= lineBuffer_2100;
    end
    if (sel) begin
      lineBuffer_2102 <= lineBuffer_2101;
    end
    if (sel) begin
      lineBuffer_2103 <= lineBuffer_2102;
    end
    if (sel) begin
      lineBuffer_2104 <= lineBuffer_2103;
    end
    if (sel) begin
      lineBuffer_2105 <= lineBuffer_2104;
    end
    if (sel) begin
      lineBuffer_2106 <= lineBuffer_2105;
    end
    if (sel) begin
      lineBuffer_2107 <= lineBuffer_2106;
    end
    if (sel) begin
      lineBuffer_2108 <= lineBuffer_2107;
    end
    if (sel) begin
      lineBuffer_2109 <= lineBuffer_2108;
    end
    if (sel) begin
      lineBuffer_2110 <= lineBuffer_2109;
    end
    if (sel) begin
      lineBuffer_2111 <= lineBuffer_2110;
    end
    if (sel) begin
      lineBuffer_2112 <= lineBuffer_2111;
    end
    if (sel) begin
      lineBuffer_2113 <= lineBuffer_2112;
    end
    if (sel) begin
      lineBuffer_2114 <= lineBuffer_2113;
    end
    if (sel) begin
      lineBuffer_2115 <= lineBuffer_2114;
    end
    if (sel) begin
      lineBuffer_2116 <= lineBuffer_2115;
    end
    if (sel) begin
      lineBuffer_2117 <= lineBuffer_2116;
    end
    if (sel) begin
      lineBuffer_2118 <= lineBuffer_2117;
    end
    if (sel) begin
      lineBuffer_2119 <= lineBuffer_2118;
    end
    if (sel) begin
      lineBuffer_2120 <= lineBuffer_2119;
    end
    if (sel) begin
      lineBuffer_2121 <= lineBuffer_2120;
    end
    if (sel) begin
      lineBuffer_2122 <= lineBuffer_2121;
    end
    if (sel) begin
      lineBuffer_2123 <= lineBuffer_2122;
    end
    if (sel) begin
      lineBuffer_2124 <= lineBuffer_2123;
    end
    if (sel) begin
      lineBuffer_2125 <= lineBuffer_2124;
    end
    if (sel) begin
      lineBuffer_2126 <= lineBuffer_2125;
    end
    if (sel) begin
      lineBuffer_2127 <= lineBuffer_2126;
    end
    if (sel) begin
      lineBuffer_2128 <= lineBuffer_2127;
    end
    if (sel) begin
      lineBuffer_2129 <= lineBuffer_2128;
    end
    if (sel) begin
      lineBuffer_2130 <= lineBuffer_2129;
    end
    if (sel) begin
      lineBuffer_2131 <= lineBuffer_2130;
    end
    if (sel) begin
      lineBuffer_2132 <= lineBuffer_2131;
    end
    if (sel) begin
      lineBuffer_2133 <= lineBuffer_2132;
    end
    if (sel) begin
      lineBuffer_2134 <= lineBuffer_2133;
    end
    if (sel) begin
      lineBuffer_2135 <= lineBuffer_2134;
    end
    if (sel) begin
      lineBuffer_2136 <= lineBuffer_2135;
    end
    if (sel) begin
      lineBuffer_2137 <= lineBuffer_2136;
    end
    if (sel) begin
      lineBuffer_2138 <= lineBuffer_2137;
    end
    if (sel) begin
      lineBuffer_2139 <= lineBuffer_2138;
    end
    if (sel) begin
      lineBuffer_2140 <= lineBuffer_2139;
    end
    if (sel) begin
      lineBuffer_2141 <= lineBuffer_2140;
    end
    if (sel) begin
      lineBuffer_2142 <= lineBuffer_2141;
    end
    if (sel) begin
      lineBuffer_2143 <= lineBuffer_2142;
    end
    if (sel) begin
      lineBuffer_2144 <= lineBuffer_2143;
    end
    if (sel) begin
      lineBuffer_2145 <= lineBuffer_2144;
    end
    if (sel) begin
      lineBuffer_2146 <= lineBuffer_2145;
    end
    if (sel) begin
      lineBuffer_2147 <= lineBuffer_2146;
    end
    if (sel) begin
      lineBuffer_2148 <= lineBuffer_2147;
    end
    if (sel) begin
      lineBuffer_2149 <= lineBuffer_2148;
    end
    if (sel) begin
      lineBuffer_2150 <= lineBuffer_2149;
    end
    if (sel) begin
      lineBuffer_2151 <= lineBuffer_2150;
    end
    if (sel) begin
      lineBuffer_2152 <= lineBuffer_2151;
    end
    if (sel) begin
      lineBuffer_2153 <= lineBuffer_2152;
    end
    if (sel) begin
      lineBuffer_2154 <= lineBuffer_2153;
    end
    if (sel) begin
      lineBuffer_2155 <= lineBuffer_2154;
    end
    if (sel) begin
      lineBuffer_2156 <= lineBuffer_2155;
    end
    if (sel) begin
      lineBuffer_2157 <= lineBuffer_2156;
    end
    if (sel) begin
      lineBuffer_2158 <= lineBuffer_2157;
    end
    if (sel) begin
      lineBuffer_2159 <= lineBuffer_2158;
    end
    if (sel) begin
      lineBuffer_2160 <= lineBuffer_2159;
    end
    if (sel) begin
      lineBuffer_2161 <= lineBuffer_2160;
    end
    if (sel) begin
      lineBuffer_2162 <= lineBuffer_2161;
    end
    if (sel) begin
      lineBuffer_2163 <= lineBuffer_2162;
    end
    if (sel) begin
      lineBuffer_2164 <= lineBuffer_2163;
    end
    if (sel) begin
      lineBuffer_2165 <= lineBuffer_2164;
    end
    if (sel) begin
      lineBuffer_2166 <= lineBuffer_2165;
    end
    if (sel) begin
      lineBuffer_2167 <= lineBuffer_2166;
    end
    if (sel) begin
      lineBuffer_2168 <= lineBuffer_2167;
    end
    if (sel) begin
      lineBuffer_2169 <= lineBuffer_2168;
    end
    if (sel) begin
      lineBuffer_2170 <= lineBuffer_2169;
    end
    if (sel) begin
      lineBuffer_2171 <= lineBuffer_2170;
    end
    if (sel) begin
      lineBuffer_2172 <= lineBuffer_2171;
    end
    if (sel) begin
      lineBuffer_2173 <= lineBuffer_2172;
    end
    if (sel) begin
      lineBuffer_2174 <= lineBuffer_2173;
    end
    if (sel) begin
      lineBuffer_2175 <= lineBuffer_2174;
    end
    if (sel) begin
      lineBuffer_2176 <= lineBuffer_2175;
    end
    if (sel) begin
      lineBuffer_2177 <= lineBuffer_2176;
    end
    if (sel) begin
      lineBuffer_2178 <= lineBuffer_2177;
    end
    if (sel) begin
      lineBuffer_2179 <= lineBuffer_2178;
    end
    if (sel) begin
      lineBuffer_2180 <= lineBuffer_2179;
    end
    if (sel) begin
      lineBuffer_2181 <= lineBuffer_2180;
    end
    if (sel) begin
      lineBuffer_2182 <= lineBuffer_2181;
    end
    if (sel) begin
      lineBuffer_2183 <= lineBuffer_2182;
    end
    if (sel) begin
      lineBuffer_2184 <= lineBuffer_2183;
    end
    if (sel) begin
      lineBuffer_2185 <= lineBuffer_2184;
    end
    if (sel) begin
      lineBuffer_2186 <= lineBuffer_2185;
    end
    if (sel) begin
      lineBuffer_2187 <= lineBuffer_2186;
    end
    if (sel) begin
      lineBuffer_2188 <= lineBuffer_2187;
    end
    if (sel) begin
      lineBuffer_2189 <= lineBuffer_2188;
    end
    if (sel) begin
      lineBuffer_2190 <= lineBuffer_2189;
    end
    if (sel) begin
      lineBuffer_2191 <= lineBuffer_2190;
    end
    if (sel) begin
      lineBuffer_2192 <= lineBuffer_2191;
    end
    if (sel) begin
      lineBuffer_2193 <= lineBuffer_2192;
    end
    if (sel) begin
      lineBuffer_2194 <= lineBuffer_2193;
    end
    if (sel) begin
      lineBuffer_2195 <= lineBuffer_2194;
    end
    if (sel) begin
      lineBuffer_2196 <= lineBuffer_2195;
    end
    if (sel) begin
      lineBuffer_2197 <= lineBuffer_2196;
    end
    if (sel) begin
      lineBuffer_2198 <= lineBuffer_2197;
    end
    if (sel) begin
      lineBuffer_2199 <= lineBuffer_2198;
    end
    if (sel) begin
      lineBuffer_2200 <= lineBuffer_2199;
    end
    if (sel) begin
      lineBuffer_2201 <= lineBuffer_2200;
    end
    if (sel) begin
      lineBuffer_2202 <= lineBuffer_2201;
    end
    if (sel) begin
      lineBuffer_2203 <= lineBuffer_2202;
    end
    if (sel) begin
      lineBuffer_2204 <= lineBuffer_2203;
    end
    if (sel) begin
      lineBuffer_2205 <= lineBuffer_2204;
    end
    if (sel) begin
      lineBuffer_2206 <= lineBuffer_2205;
    end
    if (sel) begin
      lineBuffer_2207 <= lineBuffer_2206;
    end
    if (sel) begin
      lineBuffer_2208 <= lineBuffer_2207;
    end
    if (sel) begin
      lineBuffer_2209 <= lineBuffer_2208;
    end
    if (sel) begin
      lineBuffer_2210 <= lineBuffer_2209;
    end
    if (sel) begin
      lineBuffer_2211 <= lineBuffer_2210;
    end
    if (sel) begin
      lineBuffer_2212 <= lineBuffer_2211;
    end
    if (sel) begin
      lineBuffer_2213 <= lineBuffer_2212;
    end
    if (sel) begin
      lineBuffer_2214 <= lineBuffer_2213;
    end
    if (sel) begin
      lineBuffer_2215 <= lineBuffer_2214;
    end
    if (sel) begin
      lineBuffer_2216 <= lineBuffer_2215;
    end
    if (sel) begin
      lineBuffer_2217 <= lineBuffer_2216;
    end
    if (sel) begin
      lineBuffer_2218 <= lineBuffer_2217;
    end
    if (sel) begin
      lineBuffer_2219 <= lineBuffer_2218;
    end
    if (sel) begin
      lineBuffer_2220 <= lineBuffer_2219;
    end
    if (sel) begin
      lineBuffer_2221 <= lineBuffer_2220;
    end
    if (sel) begin
      lineBuffer_2222 <= lineBuffer_2221;
    end
    if (sel) begin
      lineBuffer_2223 <= lineBuffer_2222;
    end
    if (sel) begin
      lineBuffer_2224 <= lineBuffer_2223;
    end
    if (sel) begin
      lineBuffer_2225 <= lineBuffer_2224;
    end
    if (sel) begin
      lineBuffer_2226 <= lineBuffer_2225;
    end
    if (sel) begin
      lineBuffer_2227 <= lineBuffer_2226;
    end
    if (sel) begin
      lineBuffer_2228 <= lineBuffer_2227;
    end
    if (sel) begin
      lineBuffer_2229 <= lineBuffer_2228;
    end
    if (sel) begin
      lineBuffer_2230 <= lineBuffer_2229;
    end
    if (sel) begin
      lineBuffer_2231 <= lineBuffer_2230;
    end
    if (sel) begin
      lineBuffer_2232 <= lineBuffer_2231;
    end
    if (sel) begin
      lineBuffer_2233 <= lineBuffer_2232;
    end
    if (sel) begin
      lineBuffer_2234 <= lineBuffer_2233;
    end
    if (sel) begin
      lineBuffer_2235 <= lineBuffer_2234;
    end
    if (sel) begin
      lineBuffer_2236 <= lineBuffer_2235;
    end
    if (sel) begin
      lineBuffer_2237 <= lineBuffer_2236;
    end
    if (sel) begin
      lineBuffer_2238 <= lineBuffer_2237;
    end
    if (sel) begin
      lineBuffer_2239 <= lineBuffer_2238;
    end
    if (sel) begin
      lineBuffer_2240 <= lineBuffer_2239;
    end
    if (sel) begin
      lineBuffer_2241 <= lineBuffer_2240;
    end
    if (sel) begin
      lineBuffer_2242 <= lineBuffer_2241;
    end
    if (sel) begin
      lineBuffer_2243 <= lineBuffer_2242;
    end
    if (sel) begin
      lineBuffer_2244 <= lineBuffer_2243;
    end
    if (sel) begin
      lineBuffer_2245 <= lineBuffer_2244;
    end
    if (sel) begin
      lineBuffer_2246 <= lineBuffer_2245;
    end
    if (sel) begin
      lineBuffer_2247 <= lineBuffer_2246;
    end
    if (sel) begin
      lineBuffer_2248 <= lineBuffer_2247;
    end
    if (sel) begin
      lineBuffer_2249 <= lineBuffer_2248;
    end
    if (sel) begin
      lineBuffer_2250 <= lineBuffer_2249;
    end
    if (sel) begin
      lineBuffer_2251 <= lineBuffer_2250;
    end
    if (sel) begin
      lineBuffer_2252 <= lineBuffer_2251;
    end
    if (sel) begin
      lineBuffer_2253 <= lineBuffer_2252;
    end
    if (sel) begin
      lineBuffer_2254 <= lineBuffer_2253;
    end
    if (sel) begin
      lineBuffer_2255 <= lineBuffer_2254;
    end
    if (sel) begin
      lineBuffer_2256 <= lineBuffer_2255;
    end
    if (sel) begin
      lineBuffer_2257 <= lineBuffer_2256;
    end
    if (sel) begin
      lineBuffer_2258 <= lineBuffer_2257;
    end
    if (sel) begin
      lineBuffer_2259 <= lineBuffer_2258;
    end
    if (sel) begin
      lineBuffer_2260 <= lineBuffer_2259;
    end
    if (sel) begin
      lineBuffer_2261 <= lineBuffer_2260;
    end
    if (sel) begin
      lineBuffer_2262 <= lineBuffer_2261;
    end
    if (sel) begin
      lineBuffer_2263 <= lineBuffer_2262;
    end
    if (sel) begin
      lineBuffer_2264 <= lineBuffer_2263;
    end
    if (sel) begin
      lineBuffer_2265 <= lineBuffer_2264;
    end
    if (sel) begin
      lineBuffer_2266 <= lineBuffer_2265;
    end
    if (sel) begin
      lineBuffer_2267 <= lineBuffer_2266;
    end
    if (sel) begin
      lineBuffer_2268 <= lineBuffer_2267;
    end
    if (sel) begin
      lineBuffer_2269 <= lineBuffer_2268;
    end
    if (sel) begin
      lineBuffer_2270 <= lineBuffer_2269;
    end
    if (sel) begin
      lineBuffer_2271 <= lineBuffer_2270;
    end
    if (sel) begin
      lineBuffer_2272 <= lineBuffer_2271;
    end
    if (sel) begin
      lineBuffer_2273 <= lineBuffer_2272;
    end
    if (sel) begin
      lineBuffer_2274 <= lineBuffer_2273;
    end
    if (sel) begin
      lineBuffer_2275 <= lineBuffer_2274;
    end
    if (sel) begin
      lineBuffer_2276 <= lineBuffer_2275;
    end
    if (sel) begin
      lineBuffer_2277 <= lineBuffer_2276;
    end
    if (sel) begin
      lineBuffer_2278 <= lineBuffer_2277;
    end
    if (sel) begin
      lineBuffer_2279 <= lineBuffer_2278;
    end
    if (sel) begin
      lineBuffer_2280 <= lineBuffer_2279;
    end
    if (sel) begin
      lineBuffer_2281 <= lineBuffer_2280;
    end
    if (sel) begin
      lineBuffer_2282 <= lineBuffer_2281;
    end
    if (sel) begin
      lineBuffer_2283 <= lineBuffer_2282;
    end
    if (sel) begin
      lineBuffer_2284 <= lineBuffer_2283;
    end
    if (sel) begin
      lineBuffer_2285 <= lineBuffer_2284;
    end
    if (sel) begin
      lineBuffer_2286 <= lineBuffer_2285;
    end
    if (sel) begin
      lineBuffer_2287 <= lineBuffer_2286;
    end
    if (sel) begin
      lineBuffer_2288 <= lineBuffer_2287;
    end
    if (sel) begin
      lineBuffer_2289 <= lineBuffer_2288;
    end
    if (sel) begin
      lineBuffer_2290 <= lineBuffer_2289;
    end
    if (sel) begin
      lineBuffer_2291 <= lineBuffer_2290;
    end
    if (sel) begin
      lineBuffer_2292 <= lineBuffer_2291;
    end
    if (sel) begin
      lineBuffer_2293 <= lineBuffer_2292;
    end
    if (sel) begin
      lineBuffer_2294 <= lineBuffer_2293;
    end
    if (sel) begin
      lineBuffer_2295 <= lineBuffer_2294;
    end
    if (sel) begin
      lineBuffer_2296 <= lineBuffer_2295;
    end
    if (sel) begin
      lineBuffer_2297 <= lineBuffer_2296;
    end
    if (sel) begin
      lineBuffer_2298 <= lineBuffer_2297;
    end
    if (sel) begin
      lineBuffer_2299 <= lineBuffer_2298;
    end
    if (sel) begin
      lineBuffer_2300 <= lineBuffer_2299;
    end
    if (sel) begin
      lineBuffer_2301 <= lineBuffer_2300;
    end
    if (sel) begin
      lineBuffer_2302 <= lineBuffer_2301;
    end
    if (sel) begin
      lineBuffer_2303 <= lineBuffer_2302;
    end
    if (sel) begin
      lineBuffer_2304 <= lineBuffer_2303;
    end
    if (sel) begin
      lineBuffer_2305 <= lineBuffer_2304;
    end
    if (sel) begin
      lineBuffer_2306 <= lineBuffer_2305;
    end
    if (sel) begin
      lineBuffer_2307 <= lineBuffer_2306;
    end
    if (sel) begin
      lineBuffer_2308 <= lineBuffer_2307;
    end
    if (sel) begin
      lineBuffer_2309 <= lineBuffer_2308;
    end
    if (sel) begin
      lineBuffer_2310 <= lineBuffer_2309;
    end
    if (sel) begin
      lineBuffer_2311 <= lineBuffer_2310;
    end
    if (sel) begin
      lineBuffer_2312 <= lineBuffer_2311;
    end
    if (sel) begin
      lineBuffer_2313 <= lineBuffer_2312;
    end
    if (sel) begin
      lineBuffer_2314 <= lineBuffer_2313;
    end
    if (sel) begin
      lineBuffer_2315 <= lineBuffer_2314;
    end
    if (sel) begin
      lineBuffer_2316 <= lineBuffer_2315;
    end
    if (sel) begin
      lineBuffer_2317 <= lineBuffer_2316;
    end
    if (sel) begin
      lineBuffer_2318 <= lineBuffer_2317;
    end
    if (sel) begin
      lineBuffer_2319 <= lineBuffer_2318;
    end
    if (sel) begin
      lineBuffer_2320 <= lineBuffer_2319;
    end
    if (sel) begin
      lineBuffer_2321 <= lineBuffer_2320;
    end
    if (sel) begin
      lineBuffer_2322 <= lineBuffer_2321;
    end
    if (sel) begin
      lineBuffer_2323 <= lineBuffer_2322;
    end
    if (sel) begin
      lineBuffer_2324 <= lineBuffer_2323;
    end
    if (sel) begin
      lineBuffer_2325 <= lineBuffer_2324;
    end
    if (sel) begin
      lineBuffer_2326 <= lineBuffer_2325;
    end
    if (sel) begin
      lineBuffer_2327 <= lineBuffer_2326;
    end
    if (sel) begin
      lineBuffer_2328 <= lineBuffer_2327;
    end
    if (sel) begin
      lineBuffer_2329 <= lineBuffer_2328;
    end
    if (sel) begin
      lineBuffer_2330 <= lineBuffer_2329;
    end
    if (sel) begin
      lineBuffer_2331 <= lineBuffer_2330;
    end
    if (sel) begin
      lineBuffer_2332 <= lineBuffer_2331;
    end
    if (sel) begin
      lineBuffer_2333 <= lineBuffer_2332;
    end
    if (sel) begin
      lineBuffer_2334 <= lineBuffer_2333;
    end
    if (sel) begin
      lineBuffer_2335 <= lineBuffer_2334;
    end
    if (sel) begin
      lineBuffer_2336 <= lineBuffer_2335;
    end
    if (sel) begin
      lineBuffer_2337 <= lineBuffer_2336;
    end
    if (sel) begin
      lineBuffer_2338 <= lineBuffer_2337;
    end
    if (sel) begin
      lineBuffer_2339 <= lineBuffer_2338;
    end
    if (sel) begin
      lineBuffer_2340 <= lineBuffer_2339;
    end
    if (sel) begin
      lineBuffer_2341 <= lineBuffer_2340;
    end
    if (sel) begin
      lineBuffer_2342 <= lineBuffer_2341;
    end
    if (sel) begin
      lineBuffer_2343 <= lineBuffer_2342;
    end
    if (sel) begin
      lineBuffer_2344 <= lineBuffer_2343;
    end
    if (sel) begin
      lineBuffer_2345 <= lineBuffer_2344;
    end
    if (sel) begin
      lineBuffer_2346 <= lineBuffer_2345;
    end
    if (sel) begin
      lineBuffer_2347 <= lineBuffer_2346;
    end
    if (sel) begin
      lineBuffer_2348 <= lineBuffer_2347;
    end
    if (sel) begin
      lineBuffer_2349 <= lineBuffer_2348;
    end
    if (sel) begin
      lineBuffer_2350 <= lineBuffer_2349;
    end
    if (sel) begin
      lineBuffer_2351 <= lineBuffer_2350;
    end
    if (sel) begin
      lineBuffer_2352 <= lineBuffer_2351;
    end
    if (sel) begin
      lineBuffer_2353 <= lineBuffer_2352;
    end
    if (sel) begin
      lineBuffer_2354 <= lineBuffer_2353;
    end
    if (sel) begin
      lineBuffer_2355 <= lineBuffer_2354;
    end
    if (sel) begin
      lineBuffer_2356 <= lineBuffer_2355;
    end
    if (sel) begin
      lineBuffer_2357 <= lineBuffer_2356;
    end
    if (sel) begin
      lineBuffer_2358 <= lineBuffer_2357;
    end
    if (sel) begin
      lineBuffer_2359 <= lineBuffer_2358;
    end
    if (sel) begin
      lineBuffer_2360 <= lineBuffer_2359;
    end
    if (sel) begin
      lineBuffer_2361 <= lineBuffer_2360;
    end
    if (sel) begin
      lineBuffer_2362 <= lineBuffer_2361;
    end
    if (sel) begin
      lineBuffer_2363 <= lineBuffer_2362;
    end
    if (sel) begin
      lineBuffer_2364 <= lineBuffer_2363;
    end
    if (sel) begin
      lineBuffer_2365 <= lineBuffer_2364;
    end
    if (sel) begin
      lineBuffer_2366 <= lineBuffer_2365;
    end
    if (sel) begin
      lineBuffer_2367 <= lineBuffer_2366;
    end
    if (sel) begin
      lineBuffer_2368 <= lineBuffer_2367;
    end
    if (sel) begin
      lineBuffer_2369 <= lineBuffer_2368;
    end
    if (sel) begin
      lineBuffer_2370 <= lineBuffer_2369;
    end
    if (sel) begin
      lineBuffer_2371 <= lineBuffer_2370;
    end
    if (sel) begin
      lineBuffer_2372 <= lineBuffer_2371;
    end
    if (sel) begin
      lineBuffer_2373 <= lineBuffer_2372;
    end
    if (sel) begin
      lineBuffer_2374 <= lineBuffer_2373;
    end
    if (sel) begin
      lineBuffer_2375 <= lineBuffer_2374;
    end
    if (sel) begin
      lineBuffer_2376 <= lineBuffer_2375;
    end
    if (sel) begin
      lineBuffer_2377 <= lineBuffer_2376;
    end
    if (sel) begin
      lineBuffer_2378 <= lineBuffer_2377;
    end
    if (sel) begin
      lineBuffer_2379 <= lineBuffer_2378;
    end
    if (sel) begin
      lineBuffer_2380 <= lineBuffer_2379;
    end
    if (sel) begin
      lineBuffer_2381 <= lineBuffer_2380;
    end
    if (sel) begin
      lineBuffer_2382 <= lineBuffer_2381;
    end
    if (sel) begin
      lineBuffer_2383 <= lineBuffer_2382;
    end
    if (sel) begin
      lineBuffer_2384 <= lineBuffer_2383;
    end
    if (sel) begin
      lineBuffer_2385 <= lineBuffer_2384;
    end
    if (sel) begin
      lineBuffer_2386 <= lineBuffer_2385;
    end
    if (sel) begin
      lineBuffer_2387 <= lineBuffer_2386;
    end
    if (sel) begin
      lineBuffer_2388 <= lineBuffer_2387;
    end
    if (sel) begin
      lineBuffer_2389 <= lineBuffer_2388;
    end
    if (sel) begin
      lineBuffer_2390 <= lineBuffer_2389;
    end
    if (sel) begin
      lineBuffer_2391 <= lineBuffer_2390;
    end
    if (sel) begin
      lineBuffer_2392 <= lineBuffer_2391;
    end
    if (sel) begin
      lineBuffer_2393 <= lineBuffer_2392;
    end
    if (sel) begin
      lineBuffer_2394 <= lineBuffer_2393;
    end
    if (sel) begin
      lineBuffer_2395 <= lineBuffer_2394;
    end
    if (sel) begin
      lineBuffer_2396 <= lineBuffer_2395;
    end
    if (sel) begin
      lineBuffer_2397 <= lineBuffer_2396;
    end
    if (sel) begin
      lineBuffer_2398 <= lineBuffer_2397;
    end
    if (sel) begin
      lineBuffer_2399 <= lineBuffer_2398;
    end
    if (sel) begin
      lineBuffer_2400 <= lineBuffer_2399;
    end
    if (sel) begin
      lineBuffer_2401 <= lineBuffer_2400;
    end
    if (sel) begin
      lineBuffer_2402 <= lineBuffer_2401;
    end
    if (sel) begin
      lineBuffer_2403 <= lineBuffer_2402;
    end
    if (sel) begin
      lineBuffer_2404 <= lineBuffer_2403;
    end
    if (sel) begin
      lineBuffer_2405 <= lineBuffer_2404;
    end
    if (sel) begin
      lineBuffer_2406 <= lineBuffer_2405;
    end
    if (sel) begin
      lineBuffer_2407 <= lineBuffer_2406;
    end
    if (sel) begin
      lineBuffer_2408 <= lineBuffer_2407;
    end
    if (sel) begin
      lineBuffer_2409 <= lineBuffer_2408;
    end
    if (sel) begin
      lineBuffer_2410 <= lineBuffer_2409;
    end
    if (sel) begin
      lineBuffer_2411 <= lineBuffer_2410;
    end
    if (sel) begin
      lineBuffer_2412 <= lineBuffer_2411;
    end
    if (sel) begin
      lineBuffer_2413 <= lineBuffer_2412;
    end
    if (sel) begin
      lineBuffer_2414 <= lineBuffer_2413;
    end
    if (sel) begin
      lineBuffer_2415 <= lineBuffer_2414;
    end
    if (sel) begin
      lineBuffer_2416 <= lineBuffer_2415;
    end
    if (sel) begin
      lineBuffer_2417 <= lineBuffer_2416;
    end
    if (sel) begin
      lineBuffer_2418 <= lineBuffer_2417;
    end
    if (sel) begin
      lineBuffer_2419 <= lineBuffer_2418;
    end
    if (sel) begin
      lineBuffer_2420 <= lineBuffer_2419;
    end
    if (sel) begin
      lineBuffer_2421 <= lineBuffer_2420;
    end
    if (sel) begin
      lineBuffer_2422 <= lineBuffer_2421;
    end
    if (sel) begin
      lineBuffer_2423 <= lineBuffer_2422;
    end
    if (sel) begin
      lineBuffer_2424 <= lineBuffer_2423;
    end
    if (sel) begin
      lineBuffer_2425 <= lineBuffer_2424;
    end
    if (sel) begin
      lineBuffer_2426 <= lineBuffer_2425;
    end
    if (sel) begin
      lineBuffer_2427 <= lineBuffer_2426;
    end
    if (sel) begin
      lineBuffer_2428 <= lineBuffer_2427;
    end
    if (sel) begin
      lineBuffer_2429 <= lineBuffer_2428;
    end
    if (sel) begin
      lineBuffer_2430 <= lineBuffer_2429;
    end
    if (sel) begin
      lineBuffer_2431 <= lineBuffer_2430;
    end
    if (sel) begin
      lineBuffer_2432 <= lineBuffer_2431;
    end
    if (sel) begin
      lineBuffer_2433 <= lineBuffer_2432;
    end
    if (sel) begin
      lineBuffer_2434 <= lineBuffer_2433;
    end
    if (sel) begin
      lineBuffer_2435 <= lineBuffer_2434;
    end
    if (sel) begin
      lineBuffer_2436 <= lineBuffer_2435;
    end
    if (sel) begin
      lineBuffer_2437 <= lineBuffer_2436;
    end
    if (sel) begin
      lineBuffer_2438 <= lineBuffer_2437;
    end
    if (sel) begin
      lineBuffer_2439 <= lineBuffer_2438;
    end
    if (sel) begin
      lineBuffer_2440 <= lineBuffer_2439;
    end
    if (sel) begin
      lineBuffer_2441 <= lineBuffer_2440;
    end
    if (sel) begin
      lineBuffer_2442 <= lineBuffer_2441;
    end
    if (sel) begin
      lineBuffer_2443 <= lineBuffer_2442;
    end
    if (sel) begin
      lineBuffer_2444 <= lineBuffer_2443;
    end
    if (sel) begin
      lineBuffer_2445 <= lineBuffer_2444;
    end
    if (sel) begin
      lineBuffer_2446 <= lineBuffer_2445;
    end
    if (sel) begin
      lineBuffer_2447 <= lineBuffer_2446;
    end
    if (sel) begin
      lineBuffer_2448 <= lineBuffer_2447;
    end
    if (sel) begin
      lineBuffer_2449 <= lineBuffer_2448;
    end
    if (sel) begin
      lineBuffer_2450 <= lineBuffer_2449;
    end
    if (sel) begin
      lineBuffer_2451 <= lineBuffer_2450;
    end
    if (sel) begin
      lineBuffer_2452 <= lineBuffer_2451;
    end
    if (sel) begin
      lineBuffer_2453 <= lineBuffer_2452;
    end
    if (sel) begin
      lineBuffer_2454 <= lineBuffer_2453;
    end
    if (sel) begin
      lineBuffer_2455 <= lineBuffer_2454;
    end
    if (sel) begin
      lineBuffer_2456 <= lineBuffer_2455;
    end
    if (sel) begin
      lineBuffer_2457 <= lineBuffer_2456;
    end
    if (sel) begin
      lineBuffer_2458 <= lineBuffer_2457;
    end
    if (sel) begin
      lineBuffer_2459 <= lineBuffer_2458;
    end
    if (sel) begin
      lineBuffer_2460 <= lineBuffer_2459;
    end
    if (sel) begin
      lineBuffer_2461 <= lineBuffer_2460;
    end
    if (sel) begin
      lineBuffer_2462 <= lineBuffer_2461;
    end
    if (sel) begin
      lineBuffer_2463 <= lineBuffer_2462;
    end
    if (sel) begin
      lineBuffer_2464 <= lineBuffer_2463;
    end
    if (sel) begin
      lineBuffer_2465 <= lineBuffer_2464;
    end
    if (sel) begin
      lineBuffer_2466 <= lineBuffer_2465;
    end
    if (sel) begin
      lineBuffer_2467 <= lineBuffer_2466;
    end
    if (sel) begin
      lineBuffer_2468 <= lineBuffer_2467;
    end
    if (sel) begin
      lineBuffer_2469 <= lineBuffer_2468;
    end
    if (sel) begin
      lineBuffer_2470 <= lineBuffer_2469;
    end
    if (sel) begin
      lineBuffer_2471 <= lineBuffer_2470;
    end
    if (sel) begin
      lineBuffer_2472 <= lineBuffer_2471;
    end
    if (sel) begin
      lineBuffer_2473 <= lineBuffer_2472;
    end
    if (sel) begin
      lineBuffer_2474 <= lineBuffer_2473;
    end
    if (sel) begin
      lineBuffer_2475 <= lineBuffer_2474;
    end
    if (sel) begin
      lineBuffer_2476 <= lineBuffer_2475;
    end
    if (sel) begin
      lineBuffer_2477 <= lineBuffer_2476;
    end
    if (sel) begin
      lineBuffer_2478 <= lineBuffer_2477;
    end
    if (sel) begin
      lineBuffer_2479 <= lineBuffer_2478;
    end
    if (sel) begin
      lineBuffer_2480 <= lineBuffer_2479;
    end
    if (sel) begin
      lineBuffer_2481 <= lineBuffer_2480;
    end
    if (sel) begin
      lineBuffer_2482 <= lineBuffer_2481;
    end
    if (sel) begin
      lineBuffer_2483 <= lineBuffer_2482;
    end
    if (sel) begin
      lineBuffer_2484 <= lineBuffer_2483;
    end
    if (sel) begin
      lineBuffer_2485 <= lineBuffer_2484;
    end
    if (sel) begin
      lineBuffer_2486 <= lineBuffer_2485;
    end
    if (sel) begin
      lineBuffer_2487 <= lineBuffer_2486;
    end
    if (sel) begin
      lineBuffer_2488 <= lineBuffer_2487;
    end
    if (sel) begin
      lineBuffer_2489 <= lineBuffer_2488;
    end
    if (sel) begin
      lineBuffer_2490 <= lineBuffer_2489;
    end
    if (sel) begin
      lineBuffer_2491 <= lineBuffer_2490;
    end
    if (sel) begin
      lineBuffer_2492 <= lineBuffer_2491;
    end
    if (sel) begin
      lineBuffer_2493 <= lineBuffer_2492;
    end
    if (sel) begin
      lineBuffer_2494 <= lineBuffer_2493;
    end
    if (sel) begin
      lineBuffer_2495 <= lineBuffer_2494;
    end
    if (sel) begin
      lineBuffer_2496 <= lineBuffer_2495;
    end
    if (sel) begin
      lineBuffer_2497 <= lineBuffer_2496;
    end
    if (sel) begin
      lineBuffer_2498 <= lineBuffer_2497;
    end
    if (sel) begin
      lineBuffer_2499 <= lineBuffer_2498;
    end
    if (sel) begin
      lineBuffer_2500 <= lineBuffer_2499;
    end
    if (sel) begin
      lineBuffer_2501 <= lineBuffer_2500;
    end
    if (sel) begin
      lineBuffer_2502 <= lineBuffer_2501;
    end
    if (sel) begin
      lineBuffer_2503 <= lineBuffer_2502;
    end
    if (sel) begin
      lineBuffer_2504 <= lineBuffer_2503;
    end
    if (sel) begin
      lineBuffer_2505 <= lineBuffer_2504;
    end
    if (sel) begin
      lineBuffer_2506 <= lineBuffer_2505;
    end
    if (sel) begin
      lineBuffer_2507 <= lineBuffer_2506;
    end
    if (sel) begin
      lineBuffer_2508 <= lineBuffer_2507;
    end
    if (sel) begin
      lineBuffer_2509 <= lineBuffer_2508;
    end
    if (sel) begin
      lineBuffer_2510 <= lineBuffer_2509;
    end
    if (sel) begin
      lineBuffer_2511 <= lineBuffer_2510;
    end
    if (sel) begin
      lineBuffer_2512 <= lineBuffer_2511;
    end
    if (sel) begin
      lineBuffer_2513 <= lineBuffer_2512;
    end
    if (sel) begin
      lineBuffer_2514 <= lineBuffer_2513;
    end
    if (sel) begin
      lineBuffer_2515 <= lineBuffer_2514;
    end
    if (sel) begin
      lineBuffer_2516 <= lineBuffer_2515;
    end
    if (sel) begin
      lineBuffer_2517 <= lineBuffer_2516;
    end
    if (sel) begin
      lineBuffer_2518 <= lineBuffer_2517;
    end
    if (sel) begin
      lineBuffer_2519 <= lineBuffer_2518;
    end
    if (sel) begin
      lineBuffer_2520 <= lineBuffer_2519;
    end
    if (sel) begin
      lineBuffer_2521 <= lineBuffer_2520;
    end
    if (sel) begin
      lineBuffer_2522 <= lineBuffer_2521;
    end
    if (sel) begin
      lineBuffer_2523 <= lineBuffer_2522;
    end
    if (sel) begin
      lineBuffer_2524 <= lineBuffer_2523;
    end
    if (sel) begin
      lineBuffer_2525 <= lineBuffer_2524;
    end
    if (sel) begin
      lineBuffer_2526 <= lineBuffer_2525;
    end
    if (sel) begin
      lineBuffer_2527 <= lineBuffer_2526;
    end
    if (sel) begin
      lineBuffer_2528 <= lineBuffer_2527;
    end
    if (sel) begin
      lineBuffer_2529 <= lineBuffer_2528;
    end
    if (sel) begin
      lineBuffer_2530 <= lineBuffer_2529;
    end
    if (sel) begin
      lineBuffer_2531 <= lineBuffer_2530;
    end
    if (sel) begin
      lineBuffer_2532 <= lineBuffer_2531;
    end
    if (sel) begin
      lineBuffer_2533 <= lineBuffer_2532;
    end
    if (sel) begin
      lineBuffer_2534 <= lineBuffer_2533;
    end
    if (sel) begin
      lineBuffer_2535 <= lineBuffer_2534;
    end
    if (sel) begin
      lineBuffer_2536 <= lineBuffer_2535;
    end
    if (sel) begin
      lineBuffer_2537 <= lineBuffer_2536;
    end
    if (sel) begin
      lineBuffer_2538 <= lineBuffer_2537;
    end
    if (sel) begin
      lineBuffer_2539 <= lineBuffer_2538;
    end
    if (sel) begin
      lineBuffer_2540 <= lineBuffer_2539;
    end
    if (sel) begin
      lineBuffer_2541 <= lineBuffer_2540;
    end
    if (sel) begin
      lineBuffer_2542 <= lineBuffer_2541;
    end
    if (sel) begin
      lineBuffer_2543 <= lineBuffer_2542;
    end
    if (sel) begin
      lineBuffer_2544 <= lineBuffer_2543;
    end
    if (sel) begin
      lineBuffer_2545 <= lineBuffer_2544;
    end
    if (sel) begin
      lineBuffer_2546 <= lineBuffer_2545;
    end
    if (sel) begin
      lineBuffer_2547 <= lineBuffer_2546;
    end
    if (sel) begin
      lineBuffer_2548 <= lineBuffer_2547;
    end
    if (sel) begin
      lineBuffer_2549 <= lineBuffer_2548;
    end
    if (sel) begin
      lineBuffer_2550 <= lineBuffer_2549;
    end
    if (sel) begin
      lineBuffer_2551 <= lineBuffer_2550;
    end
    if (sel) begin
      lineBuffer_2552 <= lineBuffer_2551;
    end
    if (sel) begin
      lineBuffer_2553 <= lineBuffer_2552;
    end
    if (sel) begin
      lineBuffer_2554 <= lineBuffer_2553;
    end
    if (sel) begin
      lineBuffer_2555 <= lineBuffer_2554;
    end
    if (sel) begin
      lineBuffer_2556 <= lineBuffer_2555;
    end
    if (sel) begin
      lineBuffer_2557 <= lineBuffer_2556;
    end
    if (sel) begin
      lineBuffer_2558 <= lineBuffer_2557;
    end
    if (sel) begin
      lineBuffer_2559 <= lineBuffer_2558;
    end
    if (sel) begin
      lineBuffer_2560 <= lineBuffer_2559;
    end
    if (sel) begin
      lineBuffer_2561 <= lineBuffer_2560;
    end
    if (sel) begin
      lineBuffer_2562 <= lineBuffer_2561;
    end
    if (sel) begin
      lineBuffer_2563 <= lineBuffer_2562;
    end
    if (sel) begin
      lineBuffer_2564 <= lineBuffer_2563;
    end
    if (sel) begin
      lineBuffer_2565 <= lineBuffer_2564;
    end
    if (sel) begin
      lineBuffer_2566 <= lineBuffer_2565;
    end
    if (sel) begin
      lineBuffer_2567 <= lineBuffer_2566;
    end
    if (sel) begin
      lineBuffer_2568 <= lineBuffer_2567;
    end
    if (sel) begin
      lineBuffer_2569 <= lineBuffer_2568;
    end
    if (sel) begin
      lineBuffer_2570 <= lineBuffer_2569;
    end
    if (sel) begin
      lineBuffer_2571 <= lineBuffer_2570;
    end
    if (sel) begin
      lineBuffer_2572 <= lineBuffer_2571;
    end
    if (sel) begin
      lineBuffer_2573 <= lineBuffer_2572;
    end
    if (sel) begin
      lineBuffer_2574 <= lineBuffer_2573;
    end
    if (sel) begin
      lineBuffer_2575 <= lineBuffer_2574;
    end
    if (sel) begin
      lineBuffer_2576 <= lineBuffer_2575;
    end
    if (sel) begin
      lineBuffer_2577 <= lineBuffer_2576;
    end
    if (sel) begin
      lineBuffer_2578 <= lineBuffer_2577;
    end
    if (sel) begin
      lineBuffer_2579 <= lineBuffer_2578;
    end
    if (sel) begin
      lineBuffer_2580 <= lineBuffer_2579;
    end
    if (sel) begin
      lineBuffer_2581 <= lineBuffer_2580;
    end
    if (sel) begin
      lineBuffer_2582 <= lineBuffer_2581;
    end
    if (sel) begin
      lineBuffer_2583 <= lineBuffer_2582;
    end
    if (sel) begin
      lineBuffer_2584 <= lineBuffer_2583;
    end
    if (sel) begin
      lineBuffer_2585 <= lineBuffer_2584;
    end
    if (sel) begin
      lineBuffer_2586 <= lineBuffer_2585;
    end
    if (sel) begin
      lineBuffer_2587 <= lineBuffer_2586;
    end
    if (sel) begin
      lineBuffer_2588 <= lineBuffer_2587;
    end
    if (sel) begin
      lineBuffer_2589 <= lineBuffer_2588;
    end
    if (sel) begin
      lineBuffer_2590 <= lineBuffer_2589;
    end
    if (sel) begin
      lineBuffer_2591 <= lineBuffer_2590;
    end
    if (sel) begin
      lineBuffer_2592 <= lineBuffer_2591;
    end
    if (sel) begin
      lineBuffer_2593 <= lineBuffer_2592;
    end
    if (sel) begin
      lineBuffer_2594 <= lineBuffer_2593;
    end
    if (sel) begin
      lineBuffer_2595 <= lineBuffer_2594;
    end
    if (sel) begin
      lineBuffer_2596 <= lineBuffer_2595;
    end
    if (sel) begin
      lineBuffer_2597 <= lineBuffer_2596;
    end
    if (sel) begin
      lineBuffer_2598 <= lineBuffer_2597;
    end
    if (sel) begin
      lineBuffer_2599 <= lineBuffer_2598;
    end
    if (sel) begin
      lineBuffer_2600 <= lineBuffer_2599;
    end
    if (sel) begin
      lineBuffer_2601 <= lineBuffer_2600;
    end
    if (sel) begin
      lineBuffer_2602 <= lineBuffer_2601;
    end
    if (sel) begin
      lineBuffer_2603 <= lineBuffer_2602;
    end
    if (sel) begin
      lineBuffer_2604 <= lineBuffer_2603;
    end
    if (sel) begin
      lineBuffer_2605 <= lineBuffer_2604;
    end
    if (sel) begin
      lineBuffer_2606 <= lineBuffer_2605;
    end
    if (sel) begin
      lineBuffer_2607 <= lineBuffer_2606;
    end
    if (sel) begin
      lineBuffer_2608 <= lineBuffer_2607;
    end
    if (sel) begin
      lineBuffer_2609 <= lineBuffer_2608;
    end
    if (sel) begin
      lineBuffer_2610 <= lineBuffer_2609;
    end
    if (sel) begin
      lineBuffer_2611 <= lineBuffer_2610;
    end
    if (sel) begin
      lineBuffer_2612 <= lineBuffer_2611;
    end
    if (sel) begin
      lineBuffer_2613 <= lineBuffer_2612;
    end
    if (sel) begin
      lineBuffer_2614 <= lineBuffer_2613;
    end
    if (sel) begin
      lineBuffer_2615 <= lineBuffer_2614;
    end
    if (sel) begin
      lineBuffer_2616 <= lineBuffer_2615;
    end
    if (sel) begin
      lineBuffer_2617 <= lineBuffer_2616;
    end
    if (sel) begin
      lineBuffer_2618 <= lineBuffer_2617;
    end
    if (sel) begin
      lineBuffer_2619 <= lineBuffer_2618;
    end
    if (sel) begin
      lineBuffer_2620 <= lineBuffer_2619;
    end
    if (sel) begin
      lineBuffer_2621 <= lineBuffer_2620;
    end
    if (sel) begin
      lineBuffer_2622 <= lineBuffer_2621;
    end
    if (sel) begin
      lineBuffer_2623 <= lineBuffer_2622;
    end
    if (sel) begin
      lineBuffer_2624 <= lineBuffer_2623;
    end
    if (sel) begin
      lineBuffer_2625 <= lineBuffer_2624;
    end
    if (sel) begin
      lineBuffer_2626 <= lineBuffer_2625;
    end
    if (sel) begin
      lineBuffer_2627 <= lineBuffer_2626;
    end
    if (sel) begin
      lineBuffer_2628 <= lineBuffer_2627;
    end
    if (sel) begin
      lineBuffer_2629 <= lineBuffer_2628;
    end
    if (sel) begin
      lineBuffer_2630 <= lineBuffer_2629;
    end
    if (sel) begin
      lineBuffer_2631 <= lineBuffer_2630;
    end
    if (sel) begin
      lineBuffer_2632 <= lineBuffer_2631;
    end
    if (sel) begin
      lineBuffer_2633 <= lineBuffer_2632;
    end
    if (sel) begin
      lineBuffer_2634 <= lineBuffer_2633;
    end
    if (sel) begin
      lineBuffer_2635 <= lineBuffer_2634;
    end
    if (sel) begin
      lineBuffer_2636 <= lineBuffer_2635;
    end
    if (sel) begin
      lineBuffer_2637 <= lineBuffer_2636;
    end
    if (sel) begin
      lineBuffer_2638 <= lineBuffer_2637;
    end
    if (sel) begin
      lineBuffer_2639 <= lineBuffer_2638;
    end
    if (sel) begin
      lineBuffer_2640 <= lineBuffer_2639;
    end
    if (sel) begin
      lineBuffer_2641 <= lineBuffer_2640;
    end
    if (sel) begin
      lineBuffer_2642 <= lineBuffer_2641;
    end
    if (sel) begin
      lineBuffer_2643 <= lineBuffer_2642;
    end
    if (sel) begin
      lineBuffer_2644 <= lineBuffer_2643;
    end
    if (sel) begin
      lineBuffer_2645 <= lineBuffer_2644;
    end
    if (sel) begin
      lineBuffer_2646 <= lineBuffer_2645;
    end
    if (sel) begin
      lineBuffer_2647 <= lineBuffer_2646;
    end
    if (sel) begin
      lineBuffer_2648 <= lineBuffer_2647;
    end
    if (sel) begin
      lineBuffer_2649 <= lineBuffer_2648;
    end
    if (sel) begin
      lineBuffer_2650 <= lineBuffer_2649;
    end
    if (sel) begin
      lineBuffer_2651 <= lineBuffer_2650;
    end
    if (sel) begin
      lineBuffer_2652 <= lineBuffer_2651;
    end
    if (sel) begin
      lineBuffer_2653 <= lineBuffer_2652;
    end
    if (sel) begin
      lineBuffer_2654 <= lineBuffer_2653;
    end
    if (sel) begin
      lineBuffer_2655 <= lineBuffer_2654;
    end
    if (sel) begin
      lineBuffer_2656 <= lineBuffer_2655;
    end
    if (sel) begin
      lineBuffer_2657 <= lineBuffer_2656;
    end
    if (sel) begin
      lineBuffer_2658 <= lineBuffer_2657;
    end
    if (sel) begin
      lineBuffer_2659 <= lineBuffer_2658;
    end
    if (sel) begin
      lineBuffer_2660 <= lineBuffer_2659;
    end
    if (sel) begin
      lineBuffer_2661 <= lineBuffer_2660;
    end
    if (sel) begin
      lineBuffer_2662 <= lineBuffer_2661;
    end
    if (sel) begin
      lineBuffer_2663 <= lineBuffer_2662;
    end
    if (sel) begin
      lineBuffer_2664 <= lineBuffer_2663;
    end
    if (sel) begin
      lineBuffer_2665 <= lineBuffer_2664;
    end
    if (sel) begin
      lineBuffer_2666 <= lineBuffer_2665;
    end
    if (sel) begin
      lineBuffer_2667 <= lineBuffer_2666;
    end
    if (sel) begin
      lineBuffer_2668 <= lineBuffer_2667;
    end
    if (sel) begin
      lineBuffer_2669 <= lineBuffer_2668;
    end
    if (sel) begin
      lineBuffer_2670 <= lineBuffer_2669;
    end
    if (sel) begin
      lineBuffer_2671 <= lineBuffer_2670;
    end
    if (sel) begin
      lineBuffer_2672 <= lineBuffer_2671;
    end
    if (sel) begin
      lineBuffer_2673 <= lineBuffer_2672;
    end
    if (sel) begin
      lineBuffer_2674 <= lineBuffer_2673;
    end
    if (sel) begin
      lineBuffer_2675 <= lineBuffer_2674;
    end
    if (sel) begin
      lineBuffer_2676 <= lineBuffer_2675;
    end
    if (sel) begin
      lineBuffer_2677 <= lineBuffer_2676;
    end
    if (sel) begin
      lineBuffer_2678 <= lineBuffer_2677;
    end
    if (sel) begin
      lineBuffer_2679 <= lineBuffer_2678;
    end
    if (sel) begin
      lineBuffer_2680 <= lineBuffer_2679;
    end
    if (sel) begin
      lineBuffer_2681 <= lineBuffer_2680;
    end
    if (sel) begin
      lineBuffer_2682 <= lineBuffer_2681;
    end
    if (sel) begin
      lineBuffer_2683 <= lineBuffer_2682;
    end
    if (sel) begin
      lineBuffer_2684 <= lineBuffer_2683;
    end
    if (sel) begin
      lineBuffer_2685 <= lineBuffer_2684;
    end
    if (sel) begin
      lineBuffer_2686 <= lineBuffer_2685;
    end
    if (sel) begin
      lineBuffer_2687 <= lineBuffer_2686;
    end
    if (sel) begin
      lineBuffer_2688 <= lineBuffer_2687;
    end
    if (sel) begin
      lineBuffer_2689 <= lineBuffer_2688;
    end
    if (sel) begin
      lineBuffer_2690 <= lineBuffer_2689;
    end
    if (sel) begin
      lineBuffer_2691 <= lineBuffer_2690;
    end
    if (sel) begin
      lineBuffer_2692 <= lineBuffer_2691;
    end
    if (sel) begin
      lineBuffer_2693 <= lineBuffer_2692;
    end
    if (sel) begin
      lineBuffer_2694 <= lineBuffer_2693;
    end
    if (sel) begin
      lineBuffer_2695 <= lineBuffer_2694;
    end
    if (sel) begin
      lineBuffer_2696 <= lineBuffer_2695;
    end
    if (sel) begin
      lineBuffer_2697 <= lineBuffer_2696;
    end
    if (sel) begin
      lineBuffer_2698 <= lineBuffer_2697;
    end
    if (sel) begin
      lineBuffer_2699 <= lineBuffer_2698;
    end
    if (sel) begin
      lineBuffer_2700 <= lineBuffer_2699;
    end
    if (sel) begin
      lineBuffer_2701 <= lineBuffer_2700;
    end
    if (sel) begin
      lineBuffer_2702 <= lineBuffer_2701;
    end
    if (sel) begin
      lineBuffer_2703 <= lineBuffer_2702;
    end
    if (sel) begin
      lineBuffer_2704 <= lineBuffer_2703;
    end
    if (sel) begin
      lineBuffer_2705 <= lineBuffer_2704;
    end
    if (sel) begin
      lineBuffer_2706 <= lineBuffer_2705;
    end
    if (sel) begin
      lineBuffer_2707 <= lineBuffer_2706;
    end
    if (sel) begin
      lineBuffer_2708 <= lineBuffer_2707;
    end
    if (sel) begin
      lineBuffer_2709 <= lineBuffer_2708;
    end
    if (sel) begin
      lineBuffer_2710 <= lineBuffer_2709;
    end
    if (sel) begin
      lineBuffer_2711 <= lineBuffer_2710;
    end
    if (sel) begin
      lineBuffer_2712 <= lineBuffer_2711;
    end
    if (sel) begin
      lineBuffer_2713 <= lineBuffer_2712;
    end
    if (sel) begin
      lineBuffer_2714 <= lineBuffer_2713;
    end
    if (sel) begin
      lineBuffer_2715 <= lineBuffer_2714;
    end
    if (sel) begin
      lineBuffer_2716 <= lineBuffer_2715;
    end
    if (sel) begin
      lineBuffer_2717 <= lineBuffer_2716;
    end
    if (sel) begin
      lineBuffer_2718 <= lineBuffer_2717;
    end
    if (sel) begin
      lineBuffer_2719 <= lineBuffer_2718;
    end
    if (sel) begin
      lineBuffer_2720 <= lineBuffer_2719;
    end
    if (sel) begin
      lineBuffer_2721 <= lineBuffer_2720;
    end
    if (sel) begin
      lineBuffer_2722 <= lineBuffer_2721;
    end
    if (sel) begin
      lineBuffer_2723 <= lineBuffer_2722;
    end
    if (sel) begin
      lineBuffer_2724 <= lineBuffer_2723;
    end
    if (sel) begin
      lineBuffer_2725 <= lineBuffer_2724;
    end
    if (sel) begin
      lineBuffer_2726 <= lineBuffer_2725;
    end
    if (sel) begin
      lineBuffer_2727 <= lineBuffer_2726;
    end
    if (sel) begin
      lineBuffer_2728 <= lineBuffer_2727;
    end
    if (sel) begin
      lineBuffer_2729 <= lineBuffer_2728;
    end
    if (sel) begin
      lineBuffer_2730 <= lineBuffer_2729;
    end
    if (sel) begin
      lineBuffer_2731 <= lineBuffer_2730;
    end
    if (sel) begin
      lineBuffer_2732 <= lineBuffer_2731;
    end
    if (sel) begin
      lineBuffer_2733 <= lineBuffer_2732;
    end
    if (sel) begin
      lineBuffer_2734 <= lineBuffer_2733;
    end
    if (sel) begin
      lineBuffer_2735 <= lineBuffer_2734;
    end
    if (sel) begin
      lineBuffer_2736 <= lineBuffer_2735;
    end
    if (sel) begin
      lineBuffer_2737 <= lineBuffer_2736;
    end
    if (sel) begin
      lineBuffer_2738 <= lineBuffer_2737;
    end
    if (sel) begin
      lineBuffer_2739 <= lineBuffer_2738;
    end
    if (sel) begin
      lineBuffer_2740 <= lineBuffer_2739;
    end
    if (sel) begin
      lineBuffer_2741 <= lineBuffer_2740;
    end
    if (sel) begin
      lineBuffer_2742 <= lineBuffer_2741;
    end
    if (sel) begin
      lineBuffer_2743 <= lineBuffer_2742;
    end
    if (sel) begin
      lineBuffer_2744 <= lineBuffer_2743;
    end
    if (sel) begin
      lineBuffer_2745 <= lineBuffer_2744;
    end
    if (sel) begin
      lineBuffer_2746 <= lineBuffer_2745;
    end
    if (sel) begin
      lineBuffer_2747 <= lineBuffer_2746;
    end
    if (sel) begin
      lineBuffer_2748 <= lineBuffer_2747;
    end
    if (sel) begin
      lineBuffer_2749 <= lineBuffer_2748;
    end
    if (sel) begin
      lineBuffer_2750 <= lineBuffer_2749;
    end
    if (sel) begin
      lineBuffer_2751 <= lineBuffer_2750;
    end
    if (sel) begin
      lineBuffer_2752 <= lineBuffer_2751;
    end
    if (sel) begin
      lineBuffer_2753 <= lineBuffer_2752;
    end
    if (sel) begin
      lineBuffer_2754 <= lineBuffer_2753;
    end
    if (sel) begin
      lineBuffer_2755 <= lineBuffer_2754;
    end
    if (sel) begin
      lineBuffer_2756 <= lineBuffer_2755;
    end
    if (sel) begin
      lineBuffer_2757 <= lineBuffer_2756;
    end
    if (sel) begin
      lineBuffer_2758 <= lineBuffer_2757;
    end
    if (sel) begin
      lineBuffer_2759 <= lineBuffer_2758;
    end
    if (sel) begin
      lineBuffer_2760 <= lineBuffer_2759;
    end
    if (sel) begin
      lineBuffer_2761 <= lineBuffer_2760;
    end
    if (sel) begin
      lineBuffer_2762 <= lineBuffer_2761;
    end
    if (sel) begin
      lineBuffer_2763 <= lineBuffer_2762;
    end
    if (sel) begin
      lineBuffer_2764 <= lineBuffer_2763;
    end
    if (sel) begin
      lineBuffer_2765 <= lineBuffer_2764;
    end
    if (sel) begin
      lineBuffer_2766 <= lineBuffer_2765;
    end
    if (sel) begin
      lineBuffer_2767 <= lineBuffer_2766;
    end
    if (sel) begin
      lineBuffer_2768 <= lineBuffer_2767;
    end
    if (sel) begin
      lineBuffer_2769 <= lineBuffer_2768;
    end
    if (sel) begin
      lineBuffer_2770 <= lineBuffer_2769;
    end
    if (sel) begin
      lineBuffer_2771 <= lineBuffer_2770;
    end
    if (sel) begin
      lineBuffer_2772 <= lineBuffer_2771;
    end
    if (sel) begin
      lineBuffer_2773 <= lineBuffer_2772;
    end
    if (sel) begin
      lineBuffer_2774 <= lineBuffer_2773;
    end
    if (sel) begin
      lineBuffer_2775 <= lineBuffer_2774;
    end
    if (sel) begin
      lineBuffer_2776 <= lineBuffer_2775;
    end
    if (sel) begin
      lineBuffer_2777 <= lineBuffer_2776;
    end
    if (sel) begin
      lineBuffer_2778 <= lineBuffer_2777;
    end
    if (sel) begin
      lineBuffer_2779 <= lineBuffer_2778;
    end
    if (sel) begin
      lineBuffer_2780 <= lineBuffer_2779;
    end
    if (sel) begin
      lineBuffer_2781 <= lineBuffer_2780;
    end
    if (sel) begin
      lineBuffer_2782 <= lineBuffer_2781;
    end
    if (sel) begin
      lineBuffer_2783 <= lineBuffer_2782;
    end
    if (sel) begin
      lineBuffer_2784 <= lineBuffer_2783;
    end
    if (sel) begin
      lineBuffer_2785 <= lineBuffer_2784;
    end
    if (sel) begin
      lineBuffer_2786 <= lineBuffer_2785;
    end
    if (sel) begin
      lineBuffer_2787 <= lineBuffer_2786;
    end
    if (sel) begin
      lineBuffer_2788 <= lineBuffer_2787;
    end
    if (sel) begin
      lineBuffer_2789 <= lineBuffer_2788;
    end
    if (sel) begin
      lineBuffer_2790 <= lineBuffer_2789;
    end
    if (sel) begin
      lineBuffer_2791 <= lineBuffer_2790;
    end
    if (sel) begin
      lineBuffer_2792 <= lineBuffer_2791;
    end
    if (sel) begin
      lineBuffer_2793 <= lineBuffer_2792;
    end
    if (sel) begin
      lineBuffer_2794 <= lineBuffer_2793;
    end
    if (sel) begin
      lineBuffer_2795 <= lineBuffer_2794;
    end
    if (sel) begin
      lineBuffer_2796 <= lineBuffer_2795;
    end
    if (sel) begin
      lineBuffer_2797 <= lineBuffer_2796;
    end
    if (sel) begin
      lineBuffer_2798 <= lineBuffer_2797;
    end
    if (sel) begin
      lineBuffer_2799 <= lineBuffer_2798;
    end
    if (sel) begin
      lineBuffer_2800 <= lineBuffer_2799;
    end
    if (sel) begin
      lineBuffer_2801 <= lineBuffer_2800;
    end
    if (sel) begin
      lineBuffer_2802 <= lineBuffer_2801;
    end
    if (sel) begin
      lineBuffer_2803 <= lineBuffer_2802;
    end
    if (sel) begin
      lineBuffer_2804 <= lineBuffer_2803;
    end
    if (sel) begin
      lineBuffer_2805 <= lineBuffer_2804;
    end
    if (sel) begin
      lineBuffer_2806 <= lineBuffer_2805;
    end
    if (sel) begin
      lineBuffer_2807 <= lineBuffer_2806;
    end
    if (sel) begin
      lineBuffer_2808 <= lineBuffer_2807;
    end
    if (sel) begin
      lineBuffer_2809 <= lineBuffer_2808;
    end
    if (sel) begin
      lineBuffer_2810 <= lineBuffer_2809;
    end
    if (sel) begin
      lineBuffer_2811 <= lineBuffer_2810;
    end
    if (sel) begin
      lineBuffer_2812 <= lineBuffer_2811;
    end
    if (sel) begin
      lineBuffer_2813 <= lineBuffer_2812;
    end
    if (sel) begin
      lineBuffer_2814 <= lineBuffer_2813;
    end
    if (sel) begin
      lineBuffer_2815 <= lineBuffer_2814;
    end
    if (sel) begin
      lineBuffer_2816 <= lineBuffer_2815;
    end
    if (sel) begin
      lineBuffer_2817 <= lineBuffer_2816;
    end
    if (sel) begin
      lineBuffer_2818 <= lineBuffer_2817;
    end
    if (sel) begin
      lineBuffer_2819 <= lineBuffer_2818;
    end
    if (sel) begin
      lineBuffer_2820 <= lineBuffer_2819;
    end
    if (sel) begin
      lineBuffer_2821 <= lineBuffer_2820;
    end
    if (sel) begin
      lineBuffer_2822 <= lineBuffer_2821;
    end
    if (sel) begin
      lineBuffer_2823 <= lineBuffer_2822;
    end
    if (sel) begin
      lineBuffer_2824 <= lineBuffer_2823;
    end
    if (sel) begin
      lineBuffer_2825 <= lineBuffer_2824;
    end
    if (sel) begin
      lineBuffer_2826 <= lineBuffer_2825;
    end
    if (sel) begin
      lineBuffer_2827 <= lineBuffer_2826;
    end
    if (sel) begin
      lineBuffer_2828 <= lineBuffer_2827;
    end
    if (sel) begin
      lineBuffer_2829 <= lineBuffer_2828;
    end
    if (sel) begin
      lineBuffer_2830 <= lineBuffer_2829;
    end
    if (sel) begin
      lineBuffer_2831 <= lineBuffer_2830;
    end
    if (sel) begin
      lineBuffer_2832 <= lineBuffer_2831;
    end
    if (sel) begin
      lineBuffer_2833 <= lineBuffer_2832;
    end
    if (sel) begin
      lineBuffer_2834 <= lineBuffer_2833;
    end
    if (sel) begin
      lineBuffer_2835 <= lineBuffer_2834;
    end
    if (sel) begin
      lineBuffer_2836 <= lineBuffer_2835;
    end
    if (sel) begin
      lineBuffer_2837 <= lineBuffer_2836;
    end
    if (sel) begin
      lineBuffer_2838 <= lineBuffer_2837;
    end
    if (sel) begin
      lineBuffer_2839 <= lineBuffer_2838;
    end
    if (sel) begin
      lineBuffer_2840 <= lineBuffer_2839;
    end
    if (sel) begin
      lineBuffer_2841 <= lineBuffer_2840;
    end
    if (sel) begin
      lineBuffer_2842 <= lineBuffer_2841;
    end
    if (sel) begin
      lineBuffer_2843 <= lineBuffer_2842;
    end
    if (sel) begin
      lineBuffer_2844 <= lineBuffer_2843;
    end
    if (sel) begin
      lineBuffer_2845 <= lineBuffer_2844;
    end
    if (sel) begin
      lineBuffer_2846 <= lineBuffer_2845;
    end
    if (sel) begin
      lineBuffer_2847 <= lineBuffer_2846;
    end
    if (sel) begin
      lineBuffer_2848 <= lineBuffer_2847;
    end
    if (sel) begin
      lineBuffer_2849 <= lineBuffer_2848;
    end
    if (sel) begin
      lineBuffer_2850 <= lineBuffer_2849;
    end
    if (sel) begin
      lineBuffer_2851 <= lineBuffer_2850;
    end
    if (sel) begin
      lineBuffer_2852 <= lineBuffer_2851;
    end
    if (sel) begin
      lineBuffer_2853 <= lineBuffer_2852;
    end
    if (sel) begin
      lineBuffer_2854 <= lineBuffer_2853;
    end
    if (sel) begin
      lineBuffer_2855 <= lineBuffer_2854;
    end
    if (sel) begin
      lineBuffer_2856 <= lineBuffer_2855;
    end
    if (sel) begin
      lineBuffer_2857 <= lineBuffer_2856;
    end
    if (sel) begin
      lineBuffer_2858 <= lineBuffer_2857;
    end
    if (sel) begin
      lineBuffer_2859 <= lineBuffer_2858;
    end
    if (sel) begin
      lineBuffer_2860 <= lineBuffer_2859;
    end
    if (sel) begin
      lineBuffer_2861 <= lineBuffer_2860;
    end
    if (sel) begin
      lineBuffer_2862 <= lineBuffer_2861;
    end
    if (sel) begin
      lineBuffer_2863 <= lineBuffer_2862;
    end
    if (sel) begin
      lineBuffer_2864 <= lineBuffer_2863;
    end
    if (sel) begin
      lineBuffer_2865 <= lineBuffer_2864;
    end
    if (sel) begin
      lineBuffer_2866 <= lineBuffer_2865;
    end
    if (sel) begin
      lineBuffer_2867 <= lineBuffer_2866;
    end
    if (sel) begin
      lineBuffer_2868 <= lineBuffer_2867;
    end
    if (sel) begin
      lineBuffer_2869 <= lineBuffer_2868;
    end
    if (sel) begin
      lineBuffer_2870 <= lineBuffer_2869;
    end
    if (sel) begin
      lineBuffer_2871 <= lineBuffer_2870;
    end
    if (sel) begin
      lineBuffer_2872 <= lineBuffer_2871;
    end
    if (sel) begin
      lineBuffer_2873 <= lineBuffer_2872;
    end
    if (sel) begin
      lineBuffer_2874 <= lineBuffer_2873;
    end
    if (sel) begin
      lineBuffer_2875 <= lineBuffer_2874;
    end
    if (sel) begin
      lineBuffer_2876 <= lineBuffer_2875;
    end
    if (sel) begin
      lineBuffer_2877 <= lineBuffer_2876;
    end
    if (sel) begin
      lineBuffer_2878 <= lineBuffer_2877;
    end
    if (sel) begin
      lineBuffer_2879 <= lineBuffer_2878;
    end
    if (sel) begin
      lineBuffer_2880 <= lineBuffer_2879;
    end
    if (sel) begin
      lineBuffer_2881 <= lineBuffer_2880;
    end
    if (sel) begin
      lineBuffer_2882 <= lineBuffer_2881;
    end
    if (sel) begin
      lineBuffer_2883 <= lineBuffer_2882;
    end
    if (sel) begin
      lineBuffer_2884 <= lineBuffer_2883;
    end
    if (sel) begin
      lineBuffer_2885 <= lineBuffer_2884;
    end
    if (sel) begin
      lineBuffer_2886 <= lineBuffer_2885;
    end
    if (sel) begin
      lineBuffer_2887 <= lineBuffer_2886;
    end
    if (sel) begin
      lineBuffer_2888 <= lineBuffer_2887;
    end
    if (sel) begin
      lineBuffer_2889 <= lineBuffer_2888;
    end
    if (sel) begin
      lineBuffer_2890 <= lineBuffer_2889;
    end
    if (sel) begin
      lineBuffer_2891 <= lineBuffer_2890;
    end
    if (sel) begin
      lineBuffer_2892 <= lineBuffer_2891;
    end
    if (sel) begin
      lineBuffer_2893 <= lineBuffer_2892;
    end
    if (sel) begin
      lineBuffer_2894 <= lineBuffer_2893;
    end
    if (sel) begin
      lineBuffer_2895 <= lineBuffer_2894;
    end
    if (sel) begin
      lineBuffer_2896 <= lineBuffer_2895;
    end
    if (sel) begin
      lineBuffer_2897 <= lineBuffer_2896;
    end
    if (sel) begin
      lineBuffer_2898 <= lineBuffer_2897;
    end
    if (sel) begin
      lineBuffer_2899 <= lineBuffer_2898;
    end
    if (sel) begin
      lineBuffer_2900 <= lineBuffer_2899;
    end
    if (sel) begin
      lineBuffer_2901 <= lineBuffer_2900;
    end
    if (sel) begin
      lineBuffer_2902 <= lineBuffer_2901;
    end
    if (sel) begin
      lineBuffer_2903 <= lineBuffer_2902;
    end
    if (sel) begin
      lineBuffer_2904 <= lineBuffer_2903;
    end
    if (sel) begin
      lineBuffer_2905 <= lineBuffer_2904;
    end
    if (sel) begin
      lineBuffer_2906 <= lineBuffer_2905;
    end
    if (sel) begin
      lineBuffer_2907 <= lineBuffer_2906;
    end
    if (sel) begin
      lineBuffer_2908 <= lineBuffer_2907;
    end
    if (sel) begin
      lineBuffer_2909 <= lineBuffer_2908;
    end
    if (sel) begin
      lineBuffer_2910 <= lineBuffer_2909;
    end
    if (sel) begin
      lineBuffer_2911 <= lineBuffer_2910;
    end
    if (sel) begin
      lineBuffer_2912 <= lineBuffer_2911;
    end
    if (sel) begin
      lineBuffer_2913 <= lineBuffer_2912;
    end
    if (sel) begin
      lineBuffer_2914 <= lineBuffer_2913;
    end
    if (sel) begin
      lineBuffer_2915 <= lineBuffer_2914;
    end
    if (sel) begin
      lineBuffer_2916 <= lineBuffer_2915;
    end
    if (sel) begin
      lineBuffer_2917 <= lineBuffer_2916;
    end
    if (sel) begin
      lineBuffer_2918 <= lineBuffer_2917;
    end
    if (sel) begin
      lineBuffer_2919 <= lineBuffer_2918;
    end
    if (sel) begin
      lineBuffer_2920 <= lineBuffer_2919;
    end
    if (sel) begin
      lineBuffer_2921 <= lineBuffer_2920;
    end
    if (sel) begin
      lineBuffer_2922 <= lineBuffer_2921;
    end
    if (sel) begin
      lineBuffer_2923 <= lineBuffer_2922;
    end
    if (sel) begin
      lineBuffer_2924 <= lineBuffer_2923;
    end
    if (sel) begin
      lineBuffer_2925 <= lineBuffer_2924;
    end
    if (sel) begin
      lineBuffer_2926 <= lineBuffer_2925;
    end
    if (sel) begin
      lineBuffer_2927 <= lineBuffer_2926;
    end
    if (sel) begin
      lineBuffer_2928 <= lineBuffer_2927;
    end
    if (sel) begin
      lineBuffer_2929 <= lineBuffer_2928;
    end
    if (sel) begin
      lineBuffer_2930 <= lineBuffer_2929;
    end
    if (sel) begin
      lineBuffer_2931 <= lineBuffer_2930;
    end
    if (sel) begin
      lineBuffer_2932 <= lineBuffer_2931;
    end
    if (sel) begin
      lineBuffer_2933 <= lineBuffer_2932;
    end
    if (sel) begin
      lineBuffer_2934 <= lineBuffer_2933;
    end
    if (sel) begin
      lineBuffer_2935 <= lineBuffer_2934;
    end
    if (sel) begin
      lineBuffer_2936 <= lineBuffer_2935;
    end
    if (sel) begin
      lineBuffer_2937 <= lineBuffer_2936;
    end
    if (sel) begin
      lineBuffer_2938 <= lineBuffer_2937;
    end
    if (sel) begin
      lineBuffer_2939 <= lineBuffer_2938;
    end
    if (sel) begin
      lineBuffer_2940 <= lineBuffer_2939;
    end
    if (sel) begin
      lineBuffer_2941 <= lineBuffer_2940;
    end
    if (sel) begin
      lineBuffer_2942 <= lineBuffer_2941;
    end
    if (sel) begin
      lineBuffer_2943 <= lineBuffer_2942;
    end
    if (sel) begin
      lineBuffer_2944 <= lineBuffer_2943;
    end
    if (sel) begin
      lineBuffer_2945 <= lineBuffer_2944;
    end
    if (sel) begin
      lineBuffer_2946 <= lineBuffer_2945;
    end
    if (sel) begin
      lineBuffer_2947 <= lineBuffer_2946;
    end
    if (sel) begin
      lineBuffer_2948 <= lineBuffer_2947;
    end
    if (sel) begin
      lineBuffer_2949 <= lineBuffer_2948;
    end
    if (sel) begin
      lineBuffer_2950 <= lineBuffer_2949;
    end
    if (sel) begin
      lineBuffer_2951 <= lineBuffer_2950;
    end
    if (sel) begin
      lineBuffer_2952 <= lineBuffer_2951;
    end
    if (sel) begin
      lineBuffer_2953 <= lineBuffer_2952;
    end
    if (sel) begin
      lineBuffer_2954 <= lineBuffer_2953;
    end
    if (sel) begin
      lineBuffer_2955 <= lineBuffer_2954;
    end
    if (sel) begin
      lineBuffer_2956 <= lineBuffer_2955;
    end
    if (sel) begin
      lineBuffer_2957 <= lineBuffer_2956;
    end
    if (sel) begin
      lineBuffer_2958 <= lineBuffer_2957;
    end
    if (sel) begin
      lineBuffer_2959 <= lineBuffer_2958;
    end
    if (sel) begin
      lineBuffer_2960 <= lineBuffer_2959;
    end
    if (sel) begin
      lineBuffer_2961 <= lineBuffer_2960;
    end
    if (sel) begin
      lineBuffer_2962 <= lineBuffer_2961;
    end
    if (sel) begin
      lineBuffer_2963 <= lineBuffer_2962;
    end
    if (sel) begin
      lineBuffer_2964 <= lineBuffer_2963;
    end
    if (sel) begin
      lineBuffer_2965 <= lineBuffer_2964;
    end
    if (sel) begin
      lineBuffer_2966 <= lineBuffer_2965;
    end
    if (sel) begin
      lineBuffer_2967 <= lineBuffer_2966;
    end
    if (sel) begin
      lineBuffer_2968 <= lineBuffer_2967;
    end
    if (sel) begin
      lineBuffer_2969 <= lineBuffer_2968;
    end
    if (sel) begin
      lineBuffer_2970 <= lineBuffer_2969;
    end
    if (sel) begin
      lineBuffer_2971 <= lineBuffer_2970;
    end
    if (sel) begin
      lineBuffer_2972 <= lineBuffer_2971;
    end
    if (sel) begin
      lineBuffer_2973 <= lineBuffer_2972;
    end
    if (sel) begin
      lineBuffer_2974 <= lineBuffer_2973;
    end
    if (sel) begin
      lineBuffer_2975 <= lineBuffer_2974;
    end
    if (sel) begin
      lineBuffer_2976 <= lineBuffer_2975;
    end
    if (sel) begin
      lineBuffer_2977 <= lineBuffer_2976;
    end
    if (sel) begin
      lineBuffer_2978 <= lineBuffer_2977;
    end
    if (sel) begin
      lineBuffer_2979 <= lineBuffer_2978;
    end
    if (sel) begin
      lineBuffer_2980 <= lineBuffer_2979;
    end
    if (sel) begin
      lineBuffer_2981 <= lineBuffer_2980;
    end
    if (sel) begin
      lineBuffer_2982 <= lineBuffer_2981;
    end
    if (sel) begin
      lineBuffer_2983 <= lineBuffer_2982;
    end
    if (sel) begin
      lineBuffer_2984 <= lineBuffer_2983;
    end
    if (sel) begin
      lineBuffer_2985 <= lineBuffer_2984;
    end
    if (sel) begin
      lineBuffer_2986 <= lineBuffer_2985;
    end
    if (sel) begin
      lineBuffer_2987 <= lineBuffer_2986;
    end
    if (sel) begin
      lineBuffer_2988 <= lineBuffer_2987;
    end
    if (sel) begin
      lineBuffer_2989 <= lineBuffer_2988;
    end
    if (sel) begin
      lineBuffer_2990 <= lineBuffer_2989;
    end
    if (sel) begin
      lineBuffer_2991 <= lineBuffer_2990;
    end
    if (sel) begin
      lineBuffer_2992 <= lineBuffer_2991;
    end
    if (sel) begin
      lineBuffer_2993 <= lineBuffer_2992;
    end
    if (sel) begin
      lineBuffer_2994 <= lineBuffer_2993;
    end
    if (sel) begin
      lineBuffer_2995 <= lineBuffer_2994;
    end
    if (sel) begin
      lineBuffer_2996 <= lineBuffer_2995;
    end
    if (sel) begin
      lineBuffer_2997 <= lineBuffer_2996;
    end
    if (sel) begin
      lineBuffer_2998 <= lineBuffer_2997;
    end
    if (sel) begin
      lineBuffer_2999 <= lineBuffer_2998;
    end
    if (sel) begin
      lineBuffer_3000 <= lineBuffer_2999;
    end
    if (sel) begin
      lineBuffer_3001 <= lineBuffer_3000;
    end
    if (sel) begin
      lineBuffer_3002 <= lineBuffer_3001;
    end
    if (sel) begin
      lineBuffer_3003 <= lineBuffer_3002;
    end
    if (sel) begin
      lineBuffer_3004 <= lineBuffer_3003;
    end
    if (sel) begin
      lineBuffer_3005 <= lineBuffer_3004;
    end
    if (sel) begin
      lineBuffer_3006 <= lineBuffer_3005;
    end
    if (sel) begin
      lineBuffer_3007 <= lineBuffer_3006;
    end
    if (sel) begin
      lineBuffer_3008 <= lineBuffer_3007;
    end
    if (sel) begin
      lineBuffer_3009 <= lineBuffer_3008;
    end
    if (sel) begin
      lineBuffer_3010 <= lineBuffer_3009;
    end
    if (sel) begin
      lineBuffer_3011 <= lineBuffer_3010;
    end
    if (sel) begin
      lineBuffer_3012 <= lineBuffer_3011;
    end
    if (sel) begin
      lineBuffer_3013 <= lineBuffer_3012;
    end
    if (sel) begin
      lineBuffer_3014 <= lineBuffer_3013;
    end
    if (sel) begin
      lineBuffer_3015 <= lineBuffer_3014;
    end
    if (sel) begin
      lineBuffer_3016 <= lineBuffer_3015;
    end
    if (sel) begin
      lineBuffer_3017 <= lineBuffer_3016;
    end
    if (sel) begin
      lineBuffer_3018 <= lineBuffer_3017;
    end
    if (sel) begin
      lineBuffer_3019 <= lineBuffer_3018;
    end
    if (sel) begin
      lineBuffer_3020 <= lineBuffer_3019;
    end
    if (sel) begin
      lineBuffer_3021 <= lineBuffer_3020;
    end
    if (sel) begin
      lineBuffer_3022 <= lineBuffer_3021;
    end
    if (sel) begin
      lineBuffer_3023 <= lineBuffer_3022;
    end
    if (sel) begin
      lineBuffer_3024 <= lineBuffer_3023;
    end
    if (sel) begin
      lineBuffer_3025 <= lineBuffer_3024;
    end
    if (sel) begin
      lineBuffer_3026 <= lineBuffer_3025;
    end
    if (sel) begin
      lineBuffer_3027 <= lineBuffer_3026;
    end
    if (sel) begin
      lineBuffer_3028 <= lineBuffer_3027;
    end
    if (sel) begin
      lineBuffer_3029 <= lineBuffer_3028;
    end
    if (sel) begin
      lineBuffer_3030 <= lineBuffer_3029;
    end
    if (sel) begin
      lineBuffer_3031 <= lineBuffer_3030;
    end
    if (sel) begin
      lineBuffer_3032 <= lineBuffer_3031;
    end
    if (sel) begin
      lineBuffer_3033 <= lineBuffer_3032;
    end
    if (sel) begin
      lineBuffer_3034 <= lineBuffer_3033;
    end
    if (sel) begin
      lineBuffer_3035 <= lineBuffer_3034;
    end
    if (sel) begin
      lineBuffer_3036 <= lineBuffer_3035;
    end
    if (sel) begin
      lineBuffer_3037 <= lineBuffer_3036;
    end
    if (sel) begin
      lineBuffer_3038 <= lineBuffer_3037;
    end
    if (sel) begin
      lineBuffer_3039 <= lineBuffer_3038;
    end
    if (sel) begin
      lineBuffer_3040 <= lineBuffer_3039;
    end
    if (sel) begin
      lineBuffer_3041 <= lineBuffer_3040;
    end
    if (sel) begin
      lineBuffer_3042 <= lineBuffer_3041;
    end
    if (sel) begin
      lineBuffer_3043 <= lineBuffer_3042;
    end
    if (sel) begin
      lineBuffer_3044 <= lineBuffer_3043;
    end
    if (sel) begin
      lineBuffer_3045 <= lineBuffer_3044;
    end
    if (sel) begin
      lineBuffer_3046 <= lineBuffer_3045;
    end
    if (sel) begin
      lineBuffer_3047 <= lineBuffer_3046;
    end
    if (sel) begin
      lineBuffer_3048 <= lineBuffer_3047;
    end
    if (sel) begin
      lineBuffer_3049 <= lineBuffer_3048;
    end
    if (sel) begin
      lineBuffer_3050 <= lineBuffer_3049;
    end
    if (sel) begin
      lineBuffer_3051 <= lineBuffer_3050;
    end
    if (sel) begin
      lineBuffer_3052 <= lineBuffer_3051;
    end
    if (sel) begin
      lineBuffer_3053 <= lineBuffer_3052;
    end
    if (sel) begin
      lineBuffer_3054 <= lineBuffer_3053;
    end
    if (sel) begin
      lineBuffer_3055 <= lineBuffer_3054;
    end
    if (sel) begin
      lineBuffer_3056 <= lineBuffer_3055;
    end
    if (sel) begin
      lineBuffer_3057 <= lineBuffer_3056;
    end
    if (sel) begin
      lineBuffer_3058 <= lineBuffer_3057;
    end
    if (sel) begin
      lineBuffer_3059 <= lineBuffer_3058;
    end
    if (sel) begin
      lineBuffer_3060 <= lineBuffer_3059;
    end
    if (sel) begin
      lineBuffer_3061 <= lineBuffer_3060;
    end
    if (sel) begin
      lineBuffer_3062 <= lineBuffer_3061;
    end
    if (sel) begin
      lineBuffer_3063 <= lineBuffer_3062;
    end
    if (sel) begin
      lineBuffer_3064 <= lineBuffer_3063;
    end
    if (sel) begin
      lineBuffer_3065 <= lineBuffer_3064;
    end
    if (sel) begin
      lineBuffer_3066 <= lineBuffer_3065;
    end
    if (sel) begin
      lineBuffer_3067 <= lineBuffer_3066;
    end
    if (sel) begin
      lineBuffer_3068 <= lineBuffer_3067;
    end
    if (sel) begin
      lineBuffer_3069 <= lineBuffer_3068;
    end
    if (sel) begin
      lineBuffer_3070 <= lineBuffer_3069;
    end
    if (sel) begin
      lineBuffer_3071 <= lineBuffer_3070;
    end
    if (sel) begin
      lineBuffer_3072 <= lineBuffer_3071;
    end
    if (sel) begin
      lineBuffer_3073 <= lineBuffer_3072;
    end
    if (sel) begin
      lineBuffer_3074 <= lineBuffer_3073;
    end
    if (sel) begin
      lineBuffer_3075 <= lineBuffer_3074;
    end
    if (sel) begin
      lineBuffer_3076 <= lineBuffer_3075;
    end
    if (sel) begin
      lineBuffer_3077 <= lineBuffer_3076;
    end
    if (sel) begin
      lineBuffer_3078 <= lineBuffer_3077;
    end
    if (sel) begin
      lineBuffer_3079 <= lineBuffer_3078;
    end
    if (sel) begin
      lineBuffer_3080 <= lineBuffer_3079;
    end
    if (sel) begin
      lineBuffer_3081 <= lineBuffer_3080;
    end
    if (sel) begin
      lineBuffer_3082 <= lineBuffer_3081;
    end
    if (sel) begin
      lineBuffer_3083 <= lineBuffer_3082;
    end
    if (sel) begin
      lineBuffer_3084 <= lineBuffer_3083;
    end
    if (sel) begin
      lineBuffer_3085 <= lineBuffer_3084;
    end
    if (sel) begin
      lineBuffer_3086 <= lineBuffer_3085;
    end
    if (sel) begin
      lineBuffer_3087 <= lineBuffer_3086;
    end
    if (sel) begin
      lineBuffer_3088 <= lineBuffer_3087;
    end
    if (sel) begin
      lineBuffer_3089 <= lineBuffer_3088;
    end
    if (sel) begin
      lineBuffer_3090 <= lineBuffer_3089;
    end
    if (sel) begin
      lineBuffer_3091 <= lineBuffer_3090;
    end
    if (sel) begin
      lineBuffer_3092 <= lineBuffer_3091;
    end
    if (sel) begin
      lineBuffer_3093 <= lineBuffer_3092;
    end
    if (sel) begin
      lineBuffer_3094 <= lineBuffer_3093;
    end
    if (sel) begin
      lineBuffer_3095 <= lineBuffer_3094;
    end
    if (sel) begin
      lineBuffer_3096 <= lineBuffer_3095;
    end
    if (sel) begin
      lineBuffer_3097 <= lineBuffer_3096;
    end
    if (sel) begin
      lineBuffer_3098 <= lineBuffer_3097;
    end
    if (sel) begin
      lineBuffer_3099 <= lineBuffer_3098;
    end
    if (sel) begin
      lineBuffer_3100 <= lineBuffer_3099;
    end
    if (sel) begin
      lineBuffer_3101 <= lineBuffer_3100;
    end
    if (sel) begin
      lineBuffer_3102 <= lineBuffer_3101;
    end
    if (sel) begin
      lineBuffer_3103 <= lineBuffer_3102;
    end
    if (sel) begin
      lineBuffer_3104 <= lineBuffer_3103;
    end
    if (sel) begin
      lineBuffer_3105 <= lineBuffer_3104;
    end
    if (sel) begin
      lineBuffer_3106 <= lineBuffer_3105;
    end
    if (sel) begin
      lineBuffer_3107 <= lineBuffer_3106;
    end
    if (sel) begin
      lineBuffer_3108 <= lineBuffer_3107;
    end
    if (sel) begin
      lineBuffer_3109 <= lineBuffer_3108;
    end
    if (sel) begin
      lineBuffer_3110 <= lineBuffer_3109;
    end
    if (sel) begin
      lineBuffer_3111 <= lineBuffer_3110;
    end
    if (sel) begin
      lineBuffer_3112 <= lineBuffer_3111;
    end
    if (sel) begin
      lineBuffer_3113 <= lineBuffer_3112;
    end
    if (sel) begin
      lineBuffer_3114 <= lineBuffer_3113;
    end
    if (sel) begin
      lineBuffer_3115 <= lineBuffer_3114;
    end
    if (sel) begin
      lineBuffer_3116 <= lineBuffer_3115;
    end
    if (sel) begin
      lineBuffer_3117 <= lineBuffer_3116;
    end
    if (sel) begin
      lineBuffer_3118 <= lineBuffer_3117;
    end
    if (sel) begin
      lineBuffer_3119 <= lineBuffer_3118;
    end
    if (sel) begin
      lineBuffer_3120 <= lineBuffer_3119;
    end
    if (sel) begin
      lineBuffer_3121 <= lineBuffer_3120;
    end
    if (sel) begin
      lineBuffer_3122 <= lineBuffer_3121;
    end
    if (sel) begin
      lineBuffer_3123 <= lineBuffer_3122;
    end
    if (sel) begin
      lineBuffer_3124 <= lineBuffer_3123;
    end
    if (sel) begin
      lineBuffer_3125 <= lineBuffer_3124;
    end
    if (sel) begin
      lineBuffer_3126 <= lineBuffer_3125;
    end
    if (sel) begin
      lineBuffer_3127 <= lineBuffer_3126;
    end
    if (sel) begin
      lineBuffer_3128 <= lineBuffer_3127;
    end
    if (sel) begin
      lineBuffer_3129 <= lineBuffer_3128;
    end
    if (sel) begin
      lineBuffer_3130 <= lineBuffer_3129;
    end
    if (sel) begin
      lineBuffer_3131 <= lineBuffer_3130;
    end
    if (sel) begin
      lineBuffer_3132 <= lineBuffer_3131;
    end
    if (sel) begin
      lineBuffer_3133 <= lineBuffer_3132;
    end
    if (sel) begin
      lineBuffer_3134 <= lineBuffer_3133;
    end
    if (sel) begin
      lineBuffer_3135 <= lineBuffer_3134;
    end
    if (sel) begin
      lineBuffer_3136 <= lineBuffer_3135;
    end
    if (sel) begin
      lineBuffer_3137 <= lineBuffer_3136;
    end
    if (sel) begin
      lineBuffer_3138 <= lineBuffer_3137;
    end
    if (sel) begin
      lineBuffer_3139 <= lineBuffer_3138;
    end
    if (sel) begin
      lineBuffer_3140 <= lineBuffer_3139;
    end
    if (sel) begin
      lineBuffer_3141 <= lineBuffer_3140;
    end
    if (sel) begin
      lineBuffer_3142 <= lineBuffer_3141;
    end
    if (sel) begin
      lineBuffer_3143 <= lineBuffer_3142;
    end
    if (sel) begin
      lineBuffer_3144 <= lineBuffer_3143;
    end
    if (sel) begin
      lineBuffer_3145 <= lineBuffer_3144;
    end
    if (sel) begin
      lineBuffer_3146 <= lineBuffer_3145;
    end
    if (sel) begin
      lineBuffer_3147 <= lineBuffer_3146;
    end
    if (sel) begin
      lineBuffer_3148 <= lineBuffer_3147;
    end
    if (sel) begin
      lineBuffer_3149 <= lineBuffer_3148;
    end
    if (sel) begin
      lineBuffer_3150 <= lineBuffer_3149;
    end
    if (sel) begin
      lineBuffer_3151 <= lineBuffer_3150;
    end
    if (sel) begin
      lineBuffer_3152 <= lineBuffer_3151;
    end
    if (sel) begin
      lineBuffer_3153 <= lineBuffer_3152;
    end
    if (sel) begin
      lineBuffer_3154 <= lineBuffer_3153;
    end
    if (sel) begin
      lineBuffer_3155 <= lineBuffer_3154;
    end
    if (sel) begin
      lineBuffer_3156 <= lineBuffer_3155;
    end
    if (sel) begin
      lineBuffer_3157 <= lineBuffer_3156;
    end
    if (sel) begin
      lineBuffer_3158 <= lineBuffer_3157;
    end
    if (sel) begin
      lineBuffer_3159 <= lineBuffer_3158;
    end
    if (sel) begin
      lineBuffer_3160 <= lineBuffer_3159;
    end
    if (sel) begin
      lineBuffer_3161 <= lineBuffer_3160;
    end
    if (sel) begin
      lineBuffer_3162 <= lineBuffer_3161;
    end
    if (sel) begin
      lineBuffer_3163 <= lineBuffer_3162;
    end
    if (sel) begin
      lineBuffer_3164 <= lineBuffer_3163;
    end
    if (sel) begin
      lineBuffer_3165 <= lineBuffer_3164;
    end
    if (sel) begin
      lineBuffer_3166 <= lineBuffer_3165;
    end
    if (sel) begin
      lineBuffer_3167 <= lineBuffer_3166;
    end
    if (sel) begin
      lineBuffer_3168 <= lineBuffer_3167;
    end
    if (sel) begin
      lineBuffer_3169 <= lineBuffer_3168;
    end
    if (sel) begin
      lineBuffer_3170 <= lineBuffer_3169;
    end
    if (sel) begin
      lineBuffer_3171 <= lineBuffer_3170;
    end
    if (sel) begin
      lineBuffer_3172 <= lineBuffer_3171;
    end
    if (sel) begin
      lineBuffer_3173 <= lineBuffer_3172;
    end
    if (sel) begin
      lineBuffer_3174 <= lineBuffer_3173;
    end
    if (sel) begin
      lineBuffer_3175 <= lineBuffer_3174;
    end
    if (sel) begin
      lineBuffer_3176 <= lineBuffer_3175;
    end
    if (sel) begin
      lineBuffer_3177 <= lineBuffer_3176;
    end
    if (sel) begin
      lineBuffer_3178 <= lineBuffer_3177;
    end
    if (sel) begin
      lineBuffer_3179 <= lineBuffer_3178;
    end
    if (sel) begin
      lineBuffer_3180 <= lineBuffer_3179;
    end
    if (sel) begin
      lineBuffer_3181 <= lineBuffer_3180;
    end
    if (sel) begin
      lineBuffer_3182 <= lineBuffer_3181;
    end
    if (sel) begin
      lineBuffer_3183 <= lineBuffer_3182;
    end
    if (sel) begin
      lineBuffer_3184 <= lineBuffer_3183;
    end
    if (sel) begin
      lineBuffer_3185 <= lineBuffer_3184;
    end
    if (sel) begin
      lineBuffer_3186 <= lineBuffer_3185;
    end
    if (sel) begin
      lineBuffer_3187 <= lineBuffer_3186;
    end
    if (sel) begin
      lineBuffer_3188 <= lineBuffer_3187;
    end
    if (sel) begin
      lineBuffer_3189 <= lineBuffer_3188;
    end
    if (sel) begin
      lineBuffer_3190 <= lineBuffer_3189;
    end
    if (sel) begin
      lineBuffer_3191 <= lineBuffer_3190;
    end
    if (sel) begin
      lineBuffer_3192 <= lineBuffer_3191;
    end
    if (sel) begin
      lineBuffer_3193 <= lineBuffer_3192;
    end
    if (sel) begin
      lineBuffer_3194 <= lineBuffer_3193;
    end
    if (sel) begin
      lineBuffer_3195 <= lineBuffer_3194;
    end
    if (sel) begin
      lineBuffer_3196 <= lineBuffer_3195;
    end
    if (sel) begin
      lineBuffer_3197 <= lineBuffer_3196;
    end
    if (sel) begin
      lineBuffer_3198 <= lineBuffer_3197;
    end
    if (sel) begin
      lineBuffer_3199 <= lineBuffer_3198;
    end
    if (sel) begin
      lineBuffer_3200 <= lineBuffer_3199;
    end
    if (sel) begin
      lineBuffer_3201 <= lineBuffer_3200;
    end
    if (sel) begin
      lineBuffer_3202 <= lineBuffer_3201;
    end
    if (sel) begin
      lineBuffer_3203 <= lineBuffer_3202;
    end
    if (sel) begin
      lineBuffer_3204 <= lineBuffer_3203;
    end
    if (sel) begin
      lineBuffer_3205 <= lineBuffer_3204;
    end
    if (sel) begin
      lineBuffer_3206 <= lineBuffer_3205;
    end
    if (sel) begin
      lineBuffer_3207 <= lineBuffer_3206;
    end
    if (sel) begin
      lineBuffer_3208 <= lineBuffer_3207;
    end
    if (sel) begin
      lineBuffer_3209 <= lineBuffer_3208;
    end
    if (sel) begin
      lineBuffer_3210 <= lineBuffer_3209;
    end
    if (sel) begin
      lineBuffer_3211 <= lineBuffer_3210;
    end
    if (sel) begin
      lineBuffer_3212 <= lineBuffer_3211;
    end
    if (sel) begin
      lineBuffer_3213 <= lineBuffer_3212;
    end
    if (sel) begin
      lineBuffer_3214 <= lineBuffer_3213;
    end
    if (sel) begin
      lineBuffer_3215 <= lineBuffer_3214;
    end
    if (sel) begin
      lineBuffer_3216 <= lineBuffer_3215;
    end
    if (sel) begin
      lineBuffer_3217 <= lineBuffer_3216;
    end
    if (sel) begin
      lineBuffer_3218 <= lineBuffer_3217;
    end
    if (sel) begin
      lineBuffer_3219 <= lineBuffer_3218;
    end
    if (sel) begin
      lineBuffer_3220 <= lineBuffer_3219;
    end
    if (sel) begin
      lineBuffer_3221 <= lineBuffer_3220;
    end
    if (sel) begin
      lineBuffer_3222 <= lineBuffer_3221;
    end
    if (sel) begin
      lineBuffer_3223 <= lineBuffer_3222;
    end
    if (sel) begin
      lineBuffer_3224 <= lineBuffer_3223;
    end
    if (sel) begin
      lineBuffer_3225 <= lineBuffer_3224;
    end
    if (sel) begin
      lineBuffer_3226 <= lineBuffer_3225;
    end
    if (sel) begin
      lineBuffer_3227 <= lineBuffer_3226;
    end
    if (sel) begin
      lineBuffer_3228 <= lineBuffer_3227;
    end
    if (sel) begin
      lineBuffer_3229 <= lineBuffer_3228;
    end
    if (sel) begin
      lineBuffer_3230 <= lineBuffer_3229;
    end
    if (sel) begin
      lineBuffer_3231 <= lineBuffer_3230;
    end
    if (sel) begin
      lineBuffer_3232 <= lineBuffer_3231;
    end
    if (sel) begin
      lineBuffer_3233 <= lineBuffer_3232;
    end
    if (sel) begin
      lineBuffer_3234 <= lineBuffer_3233;
    end
    if (sel) begin
      lineBuffer_3235 <= lineBuffer_3234;
    end
    if (sel) begin
      lineBuffer_3236 <= lineBuffer_3235;
    end
    if (sel) begin
      lineBuffer_3237 <= lineBuffer_3236;
    end
    if (sel) begin
      lineBuffer_3238 <= lineBuffer_3237;
    end
    if (sel) begin
      lineBuffer_3239 <= lineBuffer_3238;
    end
    if (sel) begin
      lineBuffer_3240 <= lineBuffer_3239;
    end
    if (sel) begin
      lineBuffer_3241 <= lineBuffer_3240;
    end
    if (sel) begin
      lineBuffer_3242 <= lineBuffer_3241;
    end
    if (sel) begin
      lineBuffer_3243 <= lineBuffer_3242;
    end
    if (sel) begin
      lineBuffer_3244 <= lineBuffer_3243;
    end
    if (sel) begin
      lineBuffer_3245 <= lineBuffer_3244;
    end
    if (sel) begin
      lineBuffer_3246 <= lineBuffer_3245;
    end
    if (sel) begin
      lineBuffer_3247 <= lineBuffer_3246;
    end
    if (sel) begin
      lineBuffer_3248 <= lineBuffer_3247;
    end
    if (sel) begin
      lineBuffer_3249 <= lineBuffer_3248;
    end
    if (sel) begin
      lineBuffer_3250 <= lineBuffer_3249;
    end
    if (sel) begin
      lineBuffer_3251 <= lineBuffer_3250;
    end
    if (sel) begin
      lineBuffer_3252 <= lineBuffer_3251;
    end
    if (sel) begin
      lineBuffer_3253 <= lineBuffer_3252;
    end
    if (sel) begin
      lineBuffer_3254 <= lineBuffer_3253;
    end
    if (sel) begin
      lineBuffer_3255 <= lineBuffer_3254;
    end
    if (sel) begin
      lineBuffer_3256 <= lineBuffer_3255;
    end
    if (sel) begin
      lineBuffer_3257 <= lineBuffer_3256;
    end
    if (sel) begin
      lineBuffer_3258 <= lineBuffer_3257;
    end
    if (sel) begin
      lineBuffer_3259 <= lineBuffer_3258;
    end
    if (sel) begin
      lineBuffer_3260 <= lineBuffer_3259;
    end
    if (sel) begin
      lineBuffer_3261 <= lineBuffer_3260;
    end
    if (sel) begin
      lineBuffer_3262 <= lineBuffer_3261;
    end
    if (sel) begin
      lineBuffer_3263 <= lineBuffer_3262;
    end
    if (sel) begin
      lineBuffer_3264 <= lineBuffer_3263;
    end
    if (sel) begin
      lineBuffer_3265 <= lineBuffer_3264;
    end
    if (sel) begin
      lineBuffer_3266 <= lineBuffer_3265;
    end
    if (sel) begin
      lineBuffer_3267 <= lineBuffer_3266;
    end
    if (sel) begin
      lineBuffer_3268 <= lineBuffer_3267;
    end
    if (sel) begin
      lineBuffer_3269 <= lineBuffer_3268;
    end
    if (sel) begin
      lineBuffer_3270 <= lineBuffer_3269;
    end
    if (sel) begin
      lineBuffer_3271 <= lineBuffer_3270;
    end
    if (sel) begin
      lineBuffer_3272 <= lineBuffer_3271;
    end
    if (sel) begin
      lineBuffer_3273 <= lineBuffer_3272;
    end
    if (sel) begin
      lineBuffer_3274 <= lineBuffer_3273;
    end
    if (sel) begin
      lineBuffer_3275 <= lineBuffer_3274;
    end
    if (sel) begin
      lineBuffer_3276 <= lineBuffer_3275;
    end
    if (sel) begin
      lineBuffer_3277 <= lineBuffer_3276;
    end
    if (sel) begin
      lineBuffer_3278 <= lineBuffer_3277;
    end
    if (sel) begin
      lineBuffer_3279 <= lineBuffer_3278;
    end
    if (sel) begin
      lineBuffer_3280 <= lineBuffer_3279;
    end
    if (sel) begin
      lineBuffer_3281 <= lineBuffer_3280;
    end
    if (sel) begin
      lineBuffer_3282 <= lineBuffer_3281;
    end
    if (sel) begin
      lineBuffer_3283 <= lineBuffer_3282;
    end
    if (sel) begin
      lineBuffer_3284 <= lineBuffer_3283;
    end
    if (sel) begin
      lineBuffer_3285 <= lineBuffer_3284;
    end
    if (sel) begin
      lineBuffer_3286 <= lineBuffer_3285;
    end
    if (sel) begin
      lineBuffer_3287 <= lineBuffer_3286;
    end
    if (sel) begin
      lineBuffer_3288 <= lineBuffer_3287;
    end
    if (sel) begin
      lineBuffer_3289 <= lineBuffer_3288;
    end
    if (sel) begin
      lineBuffer_3290 <= lineBuffer_3289;
    end
    if (sel) begin
      lineBuffer_3291 <= lineBuffer_3290;
    end
    if (sel) begin
      lineBuffer_3292 <= lineBuffer_3291;
    end
    if (sel) begin
      lineBuffer_3293 <= lineBuffer_3292;
    end
    if (sel) begin
      lineBuffer_3294 <= lineBuffer_3293;
    end
    if (sel) begin
      lineBuffer_3295 <= lineBuffer_3294;
    end
    if (sel) begin
      lineBuffer_3296 <= lineBuffer_3295;
    end
    if (sel) begin
      lineBuffer_3297 <= lineBuffer_3296;
    end
    if (sel) begin
      lineBuffer_3298 <= lineBuffer_3297;
    end
    if (sel) begin
      lineBuffer_3299 <= lineBuffer_3298;
    end
    if (sel) begin
      lineBuffer_3300 <= lineBuffer_3299;
    end
    if (sel) begin
      lineBuffer_3301 <= lineBuffer_3300;
    end
    if (sel) begin
      lineBuffer_3302 <= lineBuffer_3301;
    end
    if (sel) begin
      lineBuffer_3303 <= lineBuffer_3302;
    end
    if (sel) begin
      lineBuffer_3304 <= lineBuffer_3303;
    end
    if (sel) begin
      lineBuffer_3305 <= lineBuffer_3304;
    end
    if (sel) begin
      lineBuffer_3306 <= lineBuffer_3305;
    end
    if (sel) begin
      lineBuffer_3307 <= lineBuffer_3306;
    end
    if (sel) begin
      lineBuffer_3308 <= lineBuffer_3307;
    end
    if (sel) begin
      lineBuffer_3309 <= lineBuffer_3308;
    end
    if (sel) begin
      lineBuffer_3310 <= lineBuffer_3309;
    end
    if (sel) begin
      lineBuffer_3311 <= lineBuffer_3310;
    end
    if (sel) begin
      lineBuffer_3312 <= lineBuffer_3311;
    end
    if (sel) begin
      lineBuffer_3313 <= lineBuffer_3312;
    end
    if (sel) begin
      lineBuffer_3314 <= lineBuffer_3313;
    end
    if (sel) begin
      lineBuffer_3315 <= lineBuffer_3314;
    end
    if (sel) begin
      lineBuffer_3316 <= lineBuffer_3315;
    end
    if (sel) begin
      lineBuffer_3317 <= lineBuffer_3316;
    end
    if (sel) begin
      lineBuffer_3318 <= lineBuffer_3317;
    end
    if (sel) begin
      lineBuffer_3319 <= lineBuffer_3318;
    end
    if (sel) begin
      lineBuffer_3320 <= lineBuffer_3319;
    end
    if (sel) begin
      lineBuffer_3321 <= lineBuffer_3320;
    end
    if (sel) begin
      lineBuffer_3322 <= lineBuffer_3321;
    end
    if (sel) begin
      lineBuffer_3323 <= lineBuffer_3322;
    end
    if (sel) begin
      lineBuffer_3324 <= lineBuffer_3323;
    end
    if (sel) begin
      lineBuffer_3325 <= lineBuffer_3324;
    end
    if (sel) begin
      lineBuffer_3326 <= lineBuffer_3325;
    end
    if (sel) begin
      lineBuffer_3327 <= lineBuffer_3326;
    end
    if (sel) begin
      lineBuffer_3328 <= lineBuffer_3327;
    end
    if (sel) begin
      lineBuffer_3329 <= lineBuffer_3328;
    end
    if (sel) begin
      lineBuffer_3330 <= lineBuffer_3329;
    end
    if (sel) begin
      lineBuffer_3331 <= lineBuffer_3330;
    end
    if (sel) begin
      lineBuffer_3332 <= lineBuffer_3331;
    end
    if (sel) begin
      lineBuffer_3333 <= lineBuffer_3332;
    end
    if (sel) begin
      lineBuffer_3334 <= lineBuffer_3333;
    end
    if (sel) begin
      lineBuffer_3335 <= lineBuffer_3334;
    end
    if (sel) begin
      lineBuffer_3336 <= lineBuffer_3335;
    end
    if (sel) begin
      lineBuffer_3337 <= lineBuffer_3336;
    end
    if (sel) begin
      lineBuffer_3338 <= lineBuffer_3337;
    end
    if (sel) begin
      lineBuffer_3339 <= lineBuffer_3338;
    end
    if (sel) begin
      lineBuffer_3340 <= lineBuffer_3339;
    end
    if (sel) begin
      lineBuffer_3341 <= lineBuffer_3340;
    end
    if (sel) begin
      lineBuffer_3342 <= lineBuffer_3341;
    end
    if (sel) begin
      lineBuffer_3343 <= lineBuffer_3342;
    end
    if (sel) begin
      lineBuffer_3344 <= lineBuffer_3343;
    end
    if (sel) begin
      lineBuffer_3345 <= lineBuffer_3344;
    end
    if (sel) begin
      lineBuffer_3346 <= lineBuffer_3345;
    end
    if (sel) begin
      lineBuffer_3347 <= lineBuffer_3346;
    end
    if (sel) begin
      lineBuffer_3348 <= lineBuffer_3347;
    end
    if (sel) begin
      lineBuffer_3349 <= lineBuffer_3348;
    end
    if (sel) begin
      lineBuffer_3350 <= lineBuffer_3349;
    end
    if (sel) begin
      lineBuffer_3351 <= lineBuffer_3350;
    end
    if (sel) begin
      lineBuffer_3352 <= lineBuffer_3351;
    end
    if (sel) begin
      lineBuffer_3353 <= lineBuffer_3352;
    end
    if (sel) begin
      lineBuffer_3354 <= lineBuffer_3353;
    end
    if (sel) begin
      lineBuffer_3355 <= lineBuffer_3354;
    end
    if (sel) begin
      lineBuffer_3356 <= lineBuffer_3355;
    end
    if (sel) begin
      lineBuffer_3357 <= lineBuffer_3356;
    end
    if (sel) begin
      lineBuffer_3358 <= lineBuffer_3357;
    end
    if (sel) begin
      lineBuffer_3359 <= lineBuffer_3358;
    end
    if (sel) begin
      lineBuffer_3360 <= lineBuffer_3359;
    end
    if (sel) begin
      lineBuffer_3361 <= lineBuffer_3360;
    end
    if (sel) begin
      lineBuffer_3362 <= lineBuffer_3361;
    end
    if (sel) begin
      lineBuffer_3363 <= lineBuffer_3362;
    end
    if (sel) begin
      lineBuffer_3364 <= lineBuffer_3363;
    end
    if (sel) begin
      lineBuffer_3365 <= lineBuffer_3364;
    end
    if (sel) begin
      lineBuffer_3366 <= lineBuffer_3365;
    end
    if (sel) begin
      lineBuffer_3367 <= lineBuffer_3366;
    end
    if (sel) begin
      lineBuffer_3368 <= lineBuffer_3367;
    end
    if (sel) begin
      lineBuffer_3369 <= lineBuffer_3368;
    end
    if (sel) begin
      lineBuffer_3370 <= lineBuffer_3369;
    end
    if (sel) begin
      lineBuffer_3371 <= lineBuffer_3370;
    end
    if (sel) begin
      lineBuffer_3372 <= lineBuffer_3371;
    end
    if (sel) begin
      lineBuffer_3373 <= lineBuffer_3372;
    end
    if (sel) begin
      lineBuffer_3374 <= lineBuffer_3373;
    end
    if (sel) begin
      lineBuffer_3375 <= lineBuffer_3374;
    end
    if (sel) begin
      lineBuffer_3376 <= lineBuffer_3375;
    end
    if (sel) begin
      lineBuffer_3377 <= lineBuffer_3376;
    end
    if (sel) begin
      lineBuffer_3378 <= lineBuffer_3377;
    end
    if (sel) begin
      lineBuffer_3379 <= lineBuffer_3378;
    end
    if (sel) begin
      lineBuffer_3380 <= lineBuffer_3379;
    end
    if (sel) begin
      lineBuffer_3381 <= lineBuffer_3380;
    end
    if (sel) begin
      lineBuffer_3382 <= lineBuffer_3381;
    end
    if (sel) begin
      lineBuffer_3383 <= lineBuffer_3382;
    end
    if (sel) begin
      lineBuffer_3384 <= lineBuffer_3383;
    end
    if (sel) begin
      lineBuffer_3385 <= lineBuffer_3384;
    end
    if (sel) begin
      lineBuffer_3386 <= lineBuffer_3385;
    end
    if (sel) begin
      lineBuffer_3387 <= lineBuffer_3386;
    end
    if (sel) begin
      lineBuffer_3388 <= lineBuffer_3387;
    end
    if (sel) begin
      lineBuffer_3389 <= lineBuffer_3388;
    end
    if (sel) begin
      lineBuffer_3390 <= lineBuffer_3389;
    end
    if (sel) begin
      lineBuffer_3391 <= lineBuffer_3390;
    end
    if (sel) begin
      lineBuffer_3392 <= lineBuffer_3391;
    end
    if (sel) begin
      lineBuffer_3393 <= lineBuffer_3392;
    end
    if (sel) begin
      lineBuffer_3394 <= lineBuffer_3393;
    end
    if (sel) begin
      lineBuffer_3395 <= lineBuffer_3394;
    end
    if (sel) begin
      lineBuffer_3396 <= lineBuffer_3395;
    end
    if (sel) begin
      lineBuffer_3397 <= lineBuffer_3396;
    end
    if (sel) begin
      lineBuffer_3398 <= lineBuffer_3397;
    end
    if (sel) begin
      lineBuffer_3399 <= lineBuffer_3398;
    end
    if (sel) begin
      lineBuffer_3400 <= lineBuffer_3399;
    end
    if (sel) begin
      lineBuffer_3401 <= lineBuffer_3400;
    end
    if (sel) begin
      lineBuffer_3402 <= lineBuffer_3401;
    end
    if (sel) begin
      lineBuffer_3403 <= lineBuffer_3402;
    end
    if (sel) begin
      lineBuffer_3404 <= lineBuffer_3403;
    end
    if (sel) begin
      lineBuffer_3405 <= lineBuffer_3404;
    end
    if (sel) begin
      lineBuffer_3406 <= lineBuffer_3405;
    end
    if (sel) begin
      lineBuffer_3407 <= lineBuffer_3406;
    end
    if (sel) begin
      lineBuffer_3408 <= lineBuffer_3407;
    end
    if (sel) begin
      lineBuffer_3409 <= lineBuffer_3408;
    end
    if (sel) begin
      lineBuffer_3410 <= lineBuffer_3409;
    end
    if (sel) begin
      lineBuffer_3411 <= lineBuffer_3410;
    end
    if (sel) begin
      lineBuffer_3412 <= lineBuffer_3411;
    end
    if (sel) begin
      lineBuffer_3413 <= lineBuffer_3412;
    end
    if (sel) begin
      lineBuffer_3414 <= lineBuffer_3413;
    end
    if (sel) begin
      lineBuffer_3415 <= lineBuffer_3414;
    end
    if (sel) begin
      lineBuffer_3416 <= lineBuffer_3415;
    end
    if (sel) begin
      lineBuffer_3417 <= lineBuffer_3416;
    end
    if (sel) begin
      lineBuffer_3418 <= lineBuffer_3417;
    end
    if (sel) begin
      lineBuffer_3419 <= lineBuffer_3418;
    end
    if (sel) begin
      lineBuffer_3420 <= lineBuffer_3419;
    end
    if (sel) begin
      lineBuffer_3421 <= lineBuffer_3420;
    end
    if (sel) begin
      lineBuffer_3422 <= lineBuffer_3421;
    end
    if (sel) begin
      lineBuffer_3423 <= lineBuffer_3422;
    end
    if (sel) begin
      lineBuffer_3424 <= lineBuffer_3423;
    end
    if (sel) begin
      lineBuffer_3425 <= lineBuffer_3424;
    end
    if (sel) begin
      lineBuffer_3426 <= lineBuffer_3425;
    end
    if (sel) begin
      lineBuffer_3427 <= lineBuffer_3426;
    end
    if (sel) begin
      lineBuffer_3428 <= lineBuffer_3427;
    end
    if (sel) begin
      lineBuffer_3429 <= lineBuffer_3428;
    end
    if (sel) begin
      lineBuffer_3430 <= lineBuffer_3429;
    end
    if (sel) begin
      lineBuffer_3431 <= lineBuffer_3430;
    end
    if (sel) begin
      lineBuffer_3432 <= lineBuffer_3431;
    end
    if (sel) begin
      lineBuffer_3433 <= lineBuffer_3432;
    end
    if (sel) begin
      lineBuffer_3434 <= lineBuffer_3433;
    end
    if (sel) begin
      lineBuffer_3435 <= lineBuffer_3434;
    end
    if (sel) begin
      lineBuffer_3436 <= lineBuffer_3435;
    end
    if (sel) begin
      lineBuffer_3437 <= lineBuffer_3436;
    end
    if (sel) begin
      lineBuffer_3438 <= lineBuffer_3437;
    end
    if (sel) begin
      lineBuffer_3439 <= lineBuffer_3438;
    end
    if (sel) begin
      lineBuffer_3440 <= lineBuffer_3439;
    end
    if (sel) begin
      lineBuffer_3441 <= lineBuffer_3440;
    end
    if (sel) begin
      lineBuffer_3442 <= lineBuffer_3441;
    end
    if (sel) begin
      lineBuffer_3443 <= lineBuffer_3442;
    end
    if (sel) begin
      lineBuffer_3444 <= lineBuffer_3443;
    end
    if (sel) begin
      lineBuffer_3445 <= lineBuffer_3444;
    end
    if (sel) begin
      lineBuffer_3446 <= lineBuffer_3445;
    end
    if (sel) begin
      lineBuffer_3447 <= lineBuffer_3446;
    end
    if (sel) begin
      lineBuffer_3448 <= lineBuffer_3447;
    end
    if (sel) begin
      lineBuffer_3449 <= lineBuffer_3448;
    end
    if (sel) begin
      lineBuffer_3450 <= lineBuffer_3449;
    end
    if (sel) begin
      lineBuffer_3451 <= lineBuffer_3450;
    end
    if (sel) begin
      lineBuffer_3452 <= lineBuffer_3451;
    end
    if (sel) begin
      lineBuffer_3453 <= lineBuffer_3452;
    end
    if (sel) begin
      lineBuffer_3454 <= lineBuffer_3453;
    end
    if (sel) begin
      lineBuffer_3455 <= lineBuffer_3454;
    end
    if (sel) begin
      lineBuffer_3456 <= lineBuffer_3455;
    end
    if (sel) begin
      lineBuffer_3457 <= lineBuffer_3456;
    end
    if (sel) begin
      lineBuffer_3458 <= lineBuffer_3457;
    end
    if (sel) begin
      lineBuffer_3459 <= lineBuffer_3458;
    end
    if (sel) begin
      lineBuffer_3460 <= lineBuffer_3459;
    end
    if (sel) begin
      lineBuffer_3461 <= lineBuffer_3460;
    end
    if (sel) begin
      lineBuffer_3462 <= lineBuffer_3461;
    end
    if (sel) begin
      lineBuffer_3463 <= lineBuffer_3462;
    end
    if (sel) begin
      lineBuffer_3464 <= lineBuffer_3463;
    end
    if (sel) begin
      lineBuffer_3465 <= lineBuffer_3464;
    end
    if (sel) begin
      lineBuffer_3466 <= lineBuffer_3465;
    end
    if (sel) begin
      lineBuffer_3467 <= lineBuffer_3466;
    end
    if (sel) begin
      lineBuffer_3468 <= lineBuffer_3467;
    end
    if (sel) begin
      lineBuffer_3469 <= lineBuffer_3468;
    end
    if (sel) begin
      lineBuffer_3470 <= lineBuffer_3469;
    end
    if (sel) begin
      lineBuffer_3471 <= lineBuffer_3470;
    end
    if (sel) begin
      lineBuffer_3472 <= lineBuffer_3471;
    end
    if (sel) begin
      lineBuffer_3473 <= lineBuffer_3472;
    end
    if (sel) begin
      lineBuffer_3474 <= lineBuffer_3473;
    end
    if (sel) begin
      lineBuffer_3475 <= lineBuffer_3474;
    end
    if (sel) begin
      lineBuffer_3476 <= lineBuffer_3475;
    end
    if (sel) begin
      lineBuffer_3477 <= lineBuffer_3476;
    end
    if (sel) begin
      lineBuffer_3478 <= lineBuffer_3477;
    end
    if (sel) begin
      lineBuffer_3479 <= lineBuffer_3478;
    end
    if (sel) begin
      lineBuffer_3480 <= lineBuffer_3479;
    end
    if (sel) begin
      lineBuffer_3481 <= lineBuffer_3480;
    end
    if (sel) begin
      lineBuffer_3482 <= lineBuffer_3481;
    end
    if (sel) begin
      lineBuffer_3483 <= lineBuffer_3482;
    end
    if (sel) begin
      lineBuffer_3484 <= lineBuffer_3483;
    end
    if (sel) begin
      lineBuffer_3485 <= lineBuffer_3484;
    end
    if (sel) begin
      lineBuffer_3486 <= lineBuffer_3485;
    end
    if (sel) begin
      lineBuffer_3487 <= lineBuffer_3486;
    end
    if (sel) begin
      lineBuffer_3488 <= lineBuffer_3487;
    end
    if (sel) begin
      lineBuffer_3489 <= lineBuffer_3488;
    end
    if (sel) begin
      lineBuffer_3490 <= lineBuffer_3489;
    end
    if (sel) begin
      lineBuffer_3491 <= lineBuffer_3490;
    end
    if (sel) begin
      lineBuffer_3492 <= lineBuffer_3491;
    end
    if (sel) begin
      lineBuffer_3493 <= lineBuffer_3492;
    end
    if (sel) begin
      lineBuffer_3494 <= lineBuffer_3493;
    end
    if (sel) begin
      lineBuffer_3495 <= lineBuffer_3494;
    end
    if (sel) begin
      lineBuffer_3496 <= lineBuffer_3495;
    end
    if (sel) begin
      lineBuffer_3497 <= lineBuffer_3496;
    end
    if (sel) begin
      lineBuffer_3498 <= lineBuffer_3497;
    end
    if (sel) begin
      lineBuffer_3499 <= lineBuffer_3498;
    end
    if (sel) begin
      lineBuffer_3500 <= lineBuffer_3499;
    end
    if (sel) begin
      lineBuffer_3501 <= lineBuffer_3500;
    end
    if (sel) begin
      lineBuffer_3502 <= lineBuffer_3501;
    end
    if (sel) begin
      lineBuffer_3503 <= lineBuffer_3502;
    end
    if (sel) begin
      lineBuffer_3504 <= lineBuffer_3503;
    end
    if (sel) begin
      lineBuffer_3505 <= lineBuffer_3504;
    end
    if (sel) begin
      lineBuffer_3506 <= lineBuffer_3505;
    end
    if (sel) begin
      lineBuffer_3507 <= lineBuffer_3506;
    end
    if (sel) begin
      lineBuffer_3508 <= lineBuffer_3507;
    end
    if (sel) begin
      lineBuffer_3509 <= lineBuffer_3508;
    end
    if (sel) begin
      lineBuffer_3510 <= lineBuffer_3509;
    end
    if (sel) begin
      lineBuffer_3511 <= lineBuffer_3510;
    end
    if (sel) begin
      lineBuffer_3512 <= lineBuffer_3511;
    end
    if (sel) begin
      lineBuffer_3513 <= lineBuffer_3512;
    end
    if (sel) begin
      lineBuffer_3514 <= lineBuffer_3513;
    end
    if (sel) begin
      lineBuffer_3515 <= lineBuffer_3514;
    end
    if (sel) begin
      lineBuffer_3516 <= lineBuffer_3515;
    end
    if (sel) begin
      lineBuffer_3517 <= lineBuffer_3516;
    end
    if (sel) begin
      lineBuffer_3518 <= lineBuffer_3517;
    end
    if (sel) begin
      lineBuffer_3519 <= lineBuffer_3518;
    end
    if (sel) begin
      lineBuffer_3520 <= lineBuffer_3519;
    end
    if (sel) begin
      lineBuffer_3521 <= lineBuffer_3520;
    end
    if (sel) begin
      lineBuffer_3522 <= lineBuffer_3521;
    end
    if (sel) begin
      lineBuffer_3523 <= lineBuffer_3522;
    end
    if (sel) begin
      lineBuffer_3524 <= lineBuffer_3523;
    end
    if (sel) begin
      lineBuffer_3525 <= lineBuffer_3524;
    end
    if (sel) begin
      lineBuffer_3526 <= lineBuffer_3525;
    end
    if (sel) begin
      lineBuffer_3527 <= lineBuffer_3526;
    end
    if (sel) begin
      lineBuffer_3528 <= lineBuffer_3527;
    end
    if (sel) begin
      lineBuffer_3529 <= lineBuffer_3528;
    end
    if (sel) begin
      lineBuffer_3530 <= lineBuffer_3529;
    end
    if (sel) begin
      lineBuffer_3531 <= lineBuffer_3530;
    end
    if (sel) begin
      lineBuffer_3532 <= lineBuffer_3531;
    end
    if (sel) begin
      lineBuffer_3533 <= lineBuffer_3532;
    end
    if (sel) begin
      lineBuffer_3534 <= lineBuffer_3533;
    end
    if (sel) begin
      lineBuffer_3535 <= lineBuffer_3534;
    end
    if (sel) begin
      lineBuffer_3536 <= lineBuffer_3535;
    end
    if (sel) begin
      lineBuffer_3537 <= lineBuffer_3536;
    end
    if (sel) begin
      lineBuffer_3538 <= lineBuffer_3537;
    end
    if (sel) begin
      lineBuffer_3539 <= lineBuffer_3538;
    end
    if (sel) begin
      lineBuffer_3540 <= lineBuffer_3539;
    end
    if (sel) begin
      lineBuffer_3541 <= lineBuffer_3540;
    end
    if (sel) begin
      lineBuffer_3542 <= lineBuffer_3541;
    end
    if (sel) begin
      lineBuffer_3543 <= lineBuffer_3542;
    end
    if (sel) begin
      lineBuffer_3544 <= lineBuffer_3543;
    end
    if (sel) begin
      lineBuffer_3545 <= lineBuffer_3544;
    end
    if (sel) begin
      lineBuffer_3546 <= lineBuffer_3545;
    end
    if (sel) begin
      lineBuffer_3547 <= lineBuffer_3546;
    end
    if (sel) begin
      lineBuffer_3548 <= lineBuffer_3547;
    end
    if (sel) begin
      lineBuffer_3549 <= lineBuffer_3548;
    end
    if (sel) begin
      lineBuffer_3550 <= lineBuffer_3549;
    end
    if (sel) begin
      lineBuffer_3551 <= lineBuffer_3550;
    end
    if (sel) begin
      lineBuffer_3552 <= lineBuffer_3551;
    end
    if (sel) begin
      lineBuffer_3553 <= lineBuffer_3552;
    end
    if (sel) begin
      lineBuffer_3554 <= lineBuffer_3553;
    end
    if (sel) begin
      lineBuffer_3555 <= lineBuffer_3554;
    end
    if (sel) begin
      lineBuffer_3556 <= lineBuffer_3555;
    end
    if (sel) begin
      lineBuffer_3557 <= lineBuffer_3556;
    end
    if (sel) begin
      lineBuffer_3558 <= lineBuffer_3557;
    end
    if (sel) begin
      lineBuffer_3559 <= lineBuffer_3558;
    end
    if (sel) begin
      lineBuffer_3560 <= lineBuffer_3559;
    end
    if (sel) begin
      lineBuffer_3561 <= lineBuffer_3560;
    end
    if (sel) begin
      lineBuffer_3562 <= lineBuffer_3561;
    end
    if (sel) begin
      lineBuffer_3563 <= lineBuffer_3562;
    end
    if (sel) begin
      lineBuffer_3564 <= lineBuffer_3563;
    end
    if (sel) begin
      lineBuffer_3565 <= lineBuffer_3564;
    end
    if (sel) begin
      lineBuffer_3566 <= lineBuffer_3565;
    end
    if (sel) begin
      lineBuffer_3567 <= lineBuffer_3566;
    end
    if (sel) begin
      lineBuffer_3568 <= lineBuffer_3567;
    end
    if (sel) begin
      lineBuffer_3569 <= lineBuffer_3568;
    end
    if (sel) begin
      lineBuffer_3570 <= lineBuffer_3569;
    end
    if (sel) begin
      lineBuffer_3571 <= lineBuffer_3570;
    end
    if (sel) begin
      lineBuffer_3572 <= lineBuffer_3571;
    end
    if (sel) begin
      lineBuffer_3573 <= lineBuffer_3572;
    end
    if (sel) begin
      lineBuffer_3574 <= lineBuffer_3573;
    end
    if (sel) begin
      lineBuffer_3575 <= lineBuffer_3574;
    end
    if (sel) begin
      lineBuffer_3576 <= lineBuffer_3575;
    end
    if (sel) begin
      lineBuffer_3577 <= lineBuffer_3576;
    end
    if (sel) begin
      lineBuffer_3578 <= lineBuffer_3577;
    end
    if (sel) begin
      lineBuffer_3579 <= lineBuffer_3578;
    end
    if (sel) begin
      lineBuffer_3580 <= lineBuffer_3579;
    end
    if (sel) begin
      lineBuffer_3581 <= lineBuffer_3580;
    end
    if (sel) begin
      lineBuffer_3582 <= lineBuffer_3581;
    end
    if (sel) begin
      lineBuffer_3583 <= lineBuffer_3582;
    end
    if (sel) begin
      lineBuffer_3584 <= lineBuffer_3583;
    end
    if (sel) begin
      lineBuffer_3585 <= lineBuffer_3584;
    end
    if (sel) begin
      lineBuffer_3586 <= lineBuffer_3585;
    end
    if (sel) begin
      lineBuffer_3587 <= lineBuffer_3586;
    end
    if (sel) begin
      lineBuffer_3588 <= lineBuffer_3587;
    end
    if (sel) begin
      lineBuffer_3589 <= lineBuffer_3588;
    end
    if (sel) begin
      lineBuffer_3590 <= lineBuffer_3589;
    end
    if (sel) begin
      lineBuffer_3591 <= lineBuffer_3590;
    end
    if (sel) begin
      lineBuffer_3592 <= lineBuffer_3591;
    end
    if (sel) begin
      lineBuffer_3593 <= lineBuffer_3592;
    end
    if (sel) begin
      lineBuffer_3594 <= lineBuffer_3593;
    end
    if (sel) begin
      lineBuffer_3595 <= lineBuffer_3594;
    end
    if (sel) begin
      lineBuffer_3596 <= lineBuffer_3595;
    end
    if (sel) begin
      lineBuffer_3597 <= lineBuffer_3596;
    end
    if (sel) begin
      lineBuffer_3598 <= lineBuffer_3597;
    end
    if (sel) begin
      lineBuffer_3599 <= lineBuffer_3598;
    end
    if (sel) begin
      lineBuffer_3600 <= lineBuffer_3599;
    end
    if (sel) begin
      lineBuffer_3601 <= lineBuffer_3600;
    end
    if (sel) begin
      lineBuffer_3602 <= lineBuffer_3601;
    end
    if (sel) begin
      lineBuffer_3603 <= lineBuffer_3602;
    end
    if (sel) begin
      lineBuffer_3604 <= lineBuffer_3603;
    end
    if (sel) begin
      lineBuffer_3605 <= lineBuffer_3604;
    end
    if (sel) begin
      lineBuffer_3606 <= lineBuffer_3605;
    end
    if (sel) begin
      lineBuffer_3607 <= lineBuffer_3606;
    end
    if (sel) begin
      lineBuffer_3608 <= lineBuffer_3607;
    end
    if (sel) begin
      lineBuffer_3609 <= lineBuffer_3608;
    end
    if (sel) begin
      lineBuffer_3610 <= lineBuffer_3609;
    end
    if (sel) begin
      lineBuffer_3611 <= lineBuffer_3610;
    end
    if (sel) begin
      lineBuffer_3612 <= lineBuffer_3611;
    end
    if (sel) begin
      lineBuffer_3613 <= lineBuffer_3612;
    end
    if (sel) begin
      lineBuffer_3614 <= lineBuffer_3613;
    end
    if (sel) begin
      lineBuffer_3615 <= lineBuffer_3614;
    end
    if (sel) begin
      lineBuffer_3616 <= lineBuffer_3615;
    end
    if (sel) begin
      lineBuffer_3617 <= lineBuffer_3616;
    end
    if (sel) begin
      lineBuffer_3618 <= lineBuffer_3617;
    end
    if (sel) begin
      lineBuffer_3619 <= lineBuffer_3618;
    end
    if (sel) begin
      lineBuffer_3620 <= lineBuffer_3619;
    end
    if (sel) begin
      lineBuffer_3621 <= lineBuffer_3620;
    end
    if (sel) begin
      lineBuffer_3622 <= lineBuffer_3621;
    end
    if (sel) begin
      lineBuffer_3623 <= lineBuffer_3622;
    end
    if (sel) begin
      lineBuffer_3624 <= lineBuffer_3623;
    end
    if (sel) begin
      lineBuffer_3625 <= lineBuffer_3624;
    end
    if (sel) begin
      lineBuffer_3626 <= lineBuffer_3625;
    end
    if (sel) begin
      lineBuffer_3627 <= lineBuffer_3626;
    end
    if (sel) begin
      lineBuffer_3628 <= lineBuffer_3627;
    end
    if (sel) begin
      lineBuffer_3629 <= lineBuffer_3628;
    end
    if (sel) begin
      lineBuffer_3630 <= lineBuffer_3629;
    end
    if (sel) begin
      lineBuffer_3631 <= lineBuffer_3630;
    end
    if (sel) begin
      lineBuffer_3632 <= lineBuffer_3631;
    end
    if (sel) begin
      lineBuffer_3633 <= lineBuffer_3632;
    end
    if (sel) begin
      lineBuffer_3634 <= lineBuffer_3633;
    end
    if (sel) begin
      lineBuffer_3635 <= lineBuffer_3634;
    end
    if (sel) begin
      lineBuffer_3636 <= lineBuffer_3635;
    end
    if (sel) begin
      lineBuffer_3637 <= lineBuffer_3636;
    end
    if (sel) begin
      lineBuffer_3638 <= lineBuffer_3637;
    end
    if (sel) begin
      lineBuffer_3639 <= lineBuffer_3638;
    end
    if (sel) begin
      lineBuffer_3640 <= lineBuffer_3639;
    end
    if (sel) begin
      lineBuffer_3641 <= lineBuffer_3640;
    end
    if (sel) begin
      lineBuffer_3642 <= lineBuffer_3641;
    end
    if (sel) begin
      lineBuffer_3643 <= lineBuffer_3642;
    end
    if (sel) begin
      lineBuffer_3644 <= lineBuffer_3643;
    end
    if (sel) begin
      lineBuffer_3645 <= lineBuffer_3644;
    end
    if (sel) begin
      lineBuffer_3646 <= lineBuffer_3645;
    end
    if (sel) begin
      lineBuffer_3647 <= lineBuffer_3646;
    end
    if (sel) begin
      lineBuffer_3648 <= lineBuffer_3647;
    end
    if (sel) begin
      lineBuffer_3649 <= lineBuffer_3648;
    end
    if (sel) begin
      lineBuffer_3650 <= lineBuffer_3649;
    end
    if (sel) begin
      lineBuffer_3651 <= lineBuffer_3650;
    end
    if (sel) begin
      lineBuffer_3652 <= lineBuffer_3651;
    end
    if (sel) begin
      lineBuffer_3653 <= lineBuffer_3652;
    end
    if (sel) begin
      lineBuffer_3654 <= lineBuffer_3653;
    end
    if (sel) begin
      lineBuffer_3655 <= lineBuffer_3654;
    end
    if (sel) begin
      lineBuffer_3656 <= lineBuffer_3655;
    end
    if (sel) begin
      lineBuffer_3657 <= lineBuffer_3656;
    end
    if (sel) begin
      lineBuffer_3658 <= lineBuffer_3657;
    end
    if (sel) begin
      lineBuffer_3659 <= lineBuffer_3658;
    end
    if (sel) begin
      lineBuffer_3660 <= lineBuffer_3659;
    end
    if (sel) begin
      lineBuffer_3661 <= lineBuffer_3660;
    end
    if (sel) begin
      lineBuffer_3662 <= lineBuffer_3661;
    end
    if (sel) begin
      lineBuffer_3663 <= lineBuffer_3662;
    end
    if (sel) begin
      lineBuffer_3664 <= lineBuffer_3663;
    end
    if (sel) begin
      lineBuffer_3665 <= lineBuffer_3664;
    end
    if (sel) begin
      lineBuffer_3666 <= lineBuffer_3665;
    end
    if (sel) begin
      lineBuffer_3667 <= lineBuffer_3666;
    end
    if (sel) begin
      lineBuffer_3668 <= lineBuffer_3667;
    end
    if (sel) begin
      lineBuffer_3669 <= lineBuffer_3668;
    end
    if (sel) begin
      lineBuffer_3670 <= lineBuffer_3669;
    end
    if (sel) begin
      lineBuffer_3671 <= lineBuffer_3670;
    end
    if (sel) begin
      lineBuffer_3672 <= lineBuffer_3671;
    end
    if (sel) begin
      lineBuffer_3673 <= lineBuffer_3672;
    end
    if (sel) begin
      lineBuffer_3674 <= lineBuffer_3673;
    end
    if (sel) begin
      lineBuffer_3675 <= lineBuffer_3674;
    end
    if (sel) begin
      lineBuffer_3676 <= lineBuffer_3675;
    end
    if (sel) begin
      lineBuffer_3677 <= lineBuffer_3676;
    end
    if (sel) begin
      lineBuffer_3678 <= lineBuffer_3677;
    end
    if (sel) begin
      lineBuffer_3679 <= lineBuffer_3678;
    end
    if (sel) begin
      lineBuffer_3680 <= lineBuffer_3679;
    end
    if (sel) begin
      lineBuffer_3681 <= lineBuffer_3680;
    end
    if (sel) begin
      lineBuffer_3682 <= lineBuffer_3681;
    end
    if (sel) begin
      lineBuffer_3683 <= lineBuffer_3682;
    end
    if (sel) begin
      lineBuffer_3684 <= lineBuffer_3683;
    end
    if (sel) begin
      lineBuffer_3685 <= lineBuffer_3684;
    end
    if (sel) begin
      lineBuffer_3686 <= lineBuffer_3685;
    end
    if (sel) begin
      lineBuffer_3687 <= lineBuffer_3686;
    end
    if (sel) begin
      lineBuffer_3688 <= lineBuffer_3687;
    end
    if (sel) begin
      lineBuffer_3689 <= lineBuffer_3688;
    end
    if (sel) begin
      lineBuffer_3690 <= lineBuffer_3689;
    end
    if (sel) begin
      lineBuffer_3691 <= lineBuffer_3690;
    end
    if (sel) begin
      lineBuffer_3692 <= lineBuffer_3691;
    end
    if (sel) begin
      lineBuffer_3693 <= lineBuffer_3692;
    end
    if (sel) begin
      lineBuffer_3694 <= lineBuffer_3693;
    end
    if (sel) begin
      lineBuffer_3695 <= lineBuffer_3694;
    end
    if (sel) begin
      lineBuffer_3696 <= lineBuffer_3695;
    end
    if (sel) begin
      lineBuffer_3697 <= lineBuffer_3696;
    end
    if (sel) begin
      lineBuffer_3698 <= lineBuffer_3697;
    end
    if (sel) begin
      lineBuffer_3699 <= lineBuffer_3698;
    end
    if (sel) begin
      lineBuffer_3700 <= lineBuffer_3699;
    end
    if (sel) begin
      lineBuffer_3701 <= lineBuffer_3700;
    end
    if (sel) begin
      lineBuffer_3702 <= lineBuffer_3701;
    end
    if (sel) begin
      lineBuffer_3703 <= lineBuffer_3702;
    end
    if (sel) begin
      lineBuffer_3704 <= lineBuffer_3703;
    end
    if (sel) begin
      lineBuffer_3705 <= lineBuffer_3704;
    end
    if (sel) begin
      lineBuffer_3706 <= lineBuffer_3705;
    end
    if (sel) begin
      lineBuffer_3707 <= lineBuffer_3706;
    end
    if (sel) begin
      lineBuffer_3708 <= lineBuffer_3707;
    end
    if (sel) begin
      lineBuffer_3709 <= lineBuffer_3708;
    end
    if (sel) begin
      lineBuffer_3710 <= lineBuffer_3709;
    end
    if (sel) begin
      lineBuffer_3711 <= lineBuffer_3710;
    end
    if (sel) begin
      lineBuffer_3712 <= lineBuffer_3711;
    end
    if (sel) begin
      lineBuffer_3713 <= lineBuffer_3712;
    end
    if (sel) begin
      lineBuffer_3714 <= lineBuffer_3713;
    end
    if (sel) begin
      lineBuffer_3715 <= lineBuffer_3714;
    end
    if (sel) begin
      lineBuffer_3716 <= lineBuffer_3715;
    end
    if (sel) begin
      lineBuffer_3717 <= lineBuffer_3716;
    end
    if (sel) begin
      lineBuffer_3718 <= lineBuffer_3717;
    end
    if (sel) begin
      lineBuffer_3719 <= lineBuffer_3718;
    end
    if (sel) begin
      lineBuffer_3720 <= lineBuffer_3719;
    end
    if (sel) begin
      lineBuffer_3721 <= lineBuffer_3720;
    end
    if (sel) begin
      lineBuffer_3722 <= lineBuffer_3721;
    end
    if (sel) begin
      lineBuffer_3723 <= lineBuffer_3722;
    end
    if (sel) begin
      lineBuffer_3724 <= lineBuffer_3723;
    end
    if (sel) begin
      lineBuffer_3725 <= lineBuffer_3724;
    end
    if (sel) begin
      lineBuffer_3726 <= lineBuffer_3725;
    end
    if (sel) begin
      lineBuffer_3727 <= lineBuffer_3726;
    end
    if (sel) begin
      lineBuffer_3728 <= lineBuffer_3727;
    end
    if (sel) begin
      lineBuffer_3729 <= lineBuffer_3728;
    end
    if (sel) begin
      lineBuffer_3730 <= lineBuffer_3729;
    end
    if (sel) begin
      lineBuffer_3731 <= lineBuffer_3730;
    end
    if (sel) begin
      lineBuffer_3732 <= lineBuffer_3731;
    end
    if (sel) begin
      lineBuffer_3733 <= lineBuffer_3732;
    end
    if (sel) begin
      lineBuffer_3734 <= lineBuffer_3733;
    end
    if (sel) begin
      lineBuffer_3735 <= lineBuffer_3734;
    end
    if (sel) begin
      lineBuffer_3736 <= lineBuffer_3735;
    end
    if (sel) begin
      lineBuffer_3737 <= lineBuffer_3736;
    end
    if (sel) begin
      lineBuffer_3738 <= lineBuffer_3737;
    end
    if (sel) begin
      lineBuffer_3739 <= lineBuffer_3738;
    end
    if (sel) begin
      lineBuffer_3740 <= lineBuffer_3739;
    end
    if (sel) begin
      lineBuffer_3741 <= lineBuffer_3740;
    end
    if (sel) begin
      lineBuffer_3742 <= lineBuffer_3741;
    end
    if (sel) begin
      lineBuffer_3743 <= lineBuffer_3742;
    end
    if (sel) begin
      lineBuffer_3744 <= lineBuffer_3743;
    end
    if (sel) begin
      lineBuffer_3745 <= lineBuffer_3744;
    end
    if (sel) begin
      lineBuffer_3746 <= lineBuffer_3745;
    end
    if (sel) begin
      lineBuffer_3747 <= lineBuffer_3746;
    end
    if (sel) begin
      lineBuffer_3748 <= lineBuffer_3747;
    end
    if (sel) begin
      lineBuffer_3749 <= lineBuffer_3748;
    end
    if (sel) begin
      lineBuffer_3750 <= lineBuffer_3749;
    end
    if (sel) begin
      lineBuffer_3751 <= lineBuffer_3750;
    end
    if (sel) begin
      lineBuffer_3752 <= lineBuffer_3751;
    end
    if (sel) begin
      lineBuffer_3753 <= lineBuffer_3752;
    end
    if (sel) begin
      lineBuffer_3754 <= lineBuffer_3753;
    end
    if (sel) begin
      lineBuffer_3755 <= lineBuffer_3754;
    end
    if (sel) begin
      lineBuffer_3756 <= lineBuffer_3755;
    end
    if (sel) begin
      lineBuffer_3757 <= lineBuffer_3756;
    end
    if (sel) begin
      lineBuffer_3758 <= lineBuffer_3757;
    end
    if (sel) begin
      lineBuffer_3759 <= lineBuffer_3758;
    end
    if (sel) begin
      lineBuffer_3760 <= lineBuffer_3759;
    end
    if (sel) begin
      lineBuffer_3761 <= lineBuffer_3760;
    end
    if (sel) begin
      lineBuffer_3762 <= lineBuffer_3761;
    end
    if (sel) begin
      lineBuffer_3763 <= lineBuffer_3762;
    end
    if (sel) begin
      lineBuffer_3764 <= lineBuffer_3763;
    end
    if (sel) begin
      lineBuffer_3765 <= lineBuffer_3764;
    end
    if (sel) begin
      lineBuffer_3766 <= lineBuffer_3765;
    end
    if (sel) begin
      lineBuffer_3767 <= lineBuffer_3766;
    end
    if (sel) begin
      lineBuffer_3768 <= lineBuffer_3767;
    end
    if (sel) begin
      lineBuffer_3769 <= lineBuffer_3768;
    end
    if (sel) begin
      lineBuffer_3770 <= lineBuffer_3769;
    end
    if (sel) begin
      lineBuffer_3771 <= lineBuffer_3770;
    end
    if (sel) begin
      lineBuffer_3772 <= lineBuffer_3771;
    end
    if (sel) begin
      lineBuffer_3773 <= lineBuffer_3772;
    end
    if (sel) begin
      lineBuffer_3774 <= lineBuffer_3773;
    end
    if (sel) begin
      lineBuffer_3775 <= lineBuffer_3774;
    end
    if (sel) begin
      lineBuffer_3776 <= lineBuffer_3775;
    end
    if (sel) begin
      lineBuffer_3777 <= lineBuffer_3776;
    end
    if (sel) begin
      lineBuffer_3778 <= lineBuffer_3777;
    end
    if (sel) begin
      lineBuffer_3779 <= lineBuffer_3778;
    end
    if (sel) begin
      lineBuffer_3780 <= lineBuffer_3779;
    end
    if (sel) begin
      lineBuffer_3781 <= lineBuffer_3780;
    end
    if (sel) begin
      lineBuffer_3782 <= lineBuffer_3781;
    end
    if (sel) begin
      lineBuffer_3783 <= lineBuffer_3782;
    end
    if (sel) begin
      lineBuffer_3784 <= lineBuffer_3783;
    end
    if (sel) begin
      lineBuffer_3785 <= lineBuffer_3784;
    end
    if (sel) begin
      lineBuffer_3786 <= lineBuffer_3785;
    end
    if (sel) begin
      lineBuffer_3787 <= lineBuffer_3786;
    end
    if (sel) begin
      lineBuffer_3788 <= lineBuffer_3787;
    end
    if (sel) begin
      lineBuffer_3789 <= lineBuffer_3788;
    end
    if (sel) begin
      lineBuffer_3790 <= lineBuffer_3789;
    end
    if (sel) begin
      lineBuffer_3791 <= lineBuffer_3790;
    end
    if (sel) begin
      lineBuffer_3792 <= lineBuffer_3791;
    end
    if (sel) begin
      lineBuffer_3793 <= lineBuffer_3792;
    end
    if (sel) begin
      lineBuffer_3794 <= lineBuffer_3793;
    end
    if (sel) begin
      lineBuffer_3795 <= lineBuffer_3794;
    end
    if (sel) begin
      lineBuffer_3796 <= lineBuffer_3795;
    end
    if (sel) begin
      lineBuffer_3797 <= lineBuffer_3796;
    end
    if (sel) begin
      lineBuffer_3798 <= lineBuffer_3797;
    end
    if (sel) begin
      lineBuffer_3799 <= lineBuffer_3798;
    end
    if (sel) begin
      lineBuffer_3800 <= lineBuffer_3799;
    end
    if (sel) begin
      lineBuffer_3801 <= lineBuffer_3800;
    end
    if (sel) begin
      lineBuffer_3802 <= lineBuffer_3801;
    end
    if (sel) begin
      lineBuffer_3803 <= lineBuffer_3802;
    end
    if (sel) begin
      lineBuffer_3804 <= lineBuffer_3803;
    end
    if (sel) begin
      lineBuffer_3805 <= lineBuffer_3804;
    end
    if (sel) begin
      lineBuffer_3806 <= lineBuffer_3805;
    end
    if (sel) begin
      lineBuffer_3807 <= lineBuffer_3806;
    end
    if (sel) begin
      lineBuffer_3808 <= lineBuffer_3807;
    end
    if (sel) begin
      lineBuffer_3809 <= lineBuffer_3808;
    end
    if (sel) begin
      lineBuffer_3810 <= lineBuffer_3809;
    end
    if (sel) begin
      lineBuffer_3811 <= lineBuffer_3810;
    end
    if (sel) begin
      lineBuffer_3812 <= lineBuffer_3811;
    end
    if (sel) begin
      lineBuffer_3813 <= lineBuffer_3812;
    end
    if (sel) begin
      lineBuffer_3814 <= lineBuffer_3813;
    end
    if (sel) begin
      lineBuffer_3815 <= lineBuffer_3814;
    end
    if (sel) begin
      lineBuffer_3816 <= lineBuffer_3815;
    end
    if (sel) begin
      lineBuffer_3817 <= lineBuffer_3816;
    end
    if (sel) begin
      lineBuffer_3818 <= lineBuffer_3817;
    end
    if (sel) begin
      lineBuffer_3819 <= lineBuffer_3818;
    end
    if (sel) begin
      lineBuffer_3820 <= lineBuffer_3819;
    end
    if (sel) begin
      lineBuffer_3821 <= lineBuffer_3820;
    end
    if (sel) begin
      lineBuffer_3822 <= lineBuffer_3821;
    end
    if (sel) begin
      lineBuffer_3823 <= lineBuffer_3822;
    end
    if (sel) begin
      lineBuffer_3824 <= lineBuffer_3823;
    end
    if (sel) begin
      lineBuffer_3825 <= lineBuffer_3824;
    end
    if (sel) begin
      lineBuffer_3826 <= lineBuffer_3825;
    end
    if (sel) begin
      lineBuffer_3827 <= lineBuffer_3826;
    end
    if (sel) begin
      lineBuffer_3828 <= lineBuffer_3827;
    end
    if (sel) begin
      lineBuffer_3829 <= lineBuffer_3828;
    end
    if (sel) begin
      lineBuffer_3830 <= lineBuffer_3829;
    end
    if (sel) begin
      lineBuffer_3831 <= lineBuffer_3830;
    end
    if (sel) begin
      lineBuffer_3832 <= lineBuffer_3831;
    end
    if (sel) begin
      lineBuffer_3833 <= lineBuffer_3832;
    end
    if (sel) begin
      lineBuffer_3834 <= lineBuffer_3833;
    end
    if (sel) begin
      lineBuffer_3835 <= lineBuffer_3834;
    end
    if (sel) begin
      lineBuffer_3836 <= lineBuffer_3835;
    end
    if (sel) begin
      lineBuffer_3837 <= lineBuffer_3836;
    end
    if (sel) begin
      lineBuffer_3838 <= lineBuffer_3837;
    end
    if (sel) begin
      lineBuffer_3839 <= lineBuffer_3838;
    end
    if (sel) begin
      lineBuffer_3840 <= lineBuffer_3839;
    end
    if (sel) begin
      lineBuffer_3841 <= lineBuffer_3840;
    end
    if (sel) begin
      lineBuffer_3842 <= lineBuffer_3841;
    end
    if (sel) begin
      lineBuffer_3843 <= lineBuffer_3842;
    end
    if (sel) begin
      lineBuffer_3844 <= lineBuffer_3843;
    end
    if (sel) begin
      lineBuffer_3845 <= lineBuffer_3844;
    end
    if (sel) begin
      lineBuffer_3846 <= lineBuffer_3845;
    end
    if (sel) begin
      lineBuffer_3847 <= lineBuffer_3846;
    end
    if (sel) begin
      lineBuffer_3848 <= lineBuffer_3847;
    end
    if (sel) begin
      lineBuffer_3849 <= lineBuffer_3848;
    end
    if (sel) begin
      lineBuffer_3850 <= lineBuffer_3849;
    end
    if (sel) begin
      lineBuffer_3851 <= lineBuffer_3850;
    end
    if (sel) begin
      lineBuffer_3852 <= lineBuffer_3851;
    end
    if (sel) begin
      lineBuffer_3853 <= lineBuffer_3852;
    end
    if (sel) begin
      lineBuffer_3854 <= lineBuffer_3853;
    end
    if (sel) begin
      lineBuffer_3855 <= lineBuffer_3854;
    end
    if (sel) begin
      lineBuffer_3856 <= lineBuffer_3855;
    end
    if (sel) begin
      lineBuffer_3857 <= lineBuffer_3856;
    end
    if (sel) begin
      lineBuffer_3858 <= lineBuffer_3857;
    end
    if (sel) begin
      lineBuffer_3859 <= lineBuffer_3858;
    end
    if (sel) begin
      lineBuffer_3860 <= lineBuffer_3859;
    end
    if (sel) begin
      lineBuffer_3861 <= lineBuffer_3860;
    end
    if (sel) begin
      lineBuffer_3862 <= lineBuffer_3861;
    end
    if (sel) begin
      lineBuffer_3863 <= lineBuffer_3862;
    end
    if (sel) begin
      lineBuffer_3864 <= lineBuffer_3863;
    end
    if (sel) begin
      lineBuffer_3865 <= lineBuffer_3864;
    end
    if (sel) begin
      lineBuffer_3866 <= lineBuffer_3865;
    end
    if (sel) begin
      lineBuffer_3867 <= lineBuffer_3866;
    end
    if (sel) begin
      lineBuffer_3868 <= lineBuffer_3867;
    end
    if (sel) begin
      lineBuffer_3869 <= lineBuffer_3868;
    end
    if (sel) begin
      lineBuffer_3870 <= lineBuffer_3869;
    end
    if (sel) begin
      lineBuffer_3871 <= lineBuffer_3870;
    end
    if (sel) begin
      lineBuffer_3872 <= lineBuffer_3871;
    end
    if (sel) begin
      lineBuffer_3873 <= lineBuffer_3872;
    end
    if (sel) begin
      lineBuffer_3874 <= lineBuffer_3873;
    end
    if (sel) begin
      lineBuffer_3875 <= lineBuffer_3874;
    end
    if (sel) begin
      lineBuffer_3876 <= lineBuffer_3875;
    end
    if (sel) begin
      lineBuffer_3877 <= lineBuffer_3876;
    end
    if (sel) begin
      lineBuffer_3878 <= lineBuffer_3877;
    end
    if (sel) begin
      lineBuffer_3879 <= lineBuffer_3878;
    end
    if (sel) begin
      lineBuffer_3880 <= lineBuffer_3879;
    end
    if (sel) begin
      lineBuffer_3881 <= lineBuffer_3880;
    end
    if (sel) begin
      lineBuffer_3882 <= lineBuffer_3881;
    end
    if (sel) begin
      lineBuffer_3883 <= lineBuffer_3882;
    end
    if (sel) begin
      lineBuffer_3884 <= lineBuffer_3883;
    end
    if (sel) begin
      lineBuffer_3885 <= lineBuffer_3884;
    end
    if (sel) begin
      lineBuffer_3886 <= lineBuffer_3885;
    end
    if (sel) begin
      lineBuffer_3887 <= lineBuffer_3886;
    end
    if (sel) begin
      lineBuffer_3888 <= lineBuffer_3887;
    end
    if (sel) begin
      lineBuffer_3889 <= lineBuffer_3888;
    end
    if (sel) begin
      lineBuffer_3890 <= lineBuffer_3889;
    end
    if (sel) begin
      lineBuffer_3891 <= lineBuffer_3890;
    end
    if (sel) begin
      lineBuffer_3892 <= lineBuffer_3891;
    end
    if (sel) begin
      lineBuffer_3893 <= lineBuffer_3892;
    end
    if (sel) begin
      lineBuffer_3894 <= lineBuffer_3893;
    end
    if (sel) begin
      lineBuffer_3895 <= lineBuffer_3894;
    end
    if (sel) begin
      lineBuffer_3896 <= lineBuffer_3895;
    end
    if (sel) begin
      lineBuffer_3897 <= lineBuffer_3896;
    end
    if (sel) begin
      lineBuffer_3898 <= lineBuffer_3897;
    end
    if (sel) begin
      lineBuffer_3899 <= lineBuffer_3898;
    end
    if (sel) begin
      lineBuffer_3900 <= lineBuffer_3899;
    end
    if (sel) begin
      lineBuffer_3901 <= lineBuffer_3900;
    end
    if (sel) begin
      lineBuffer_3902 <= lineBuffer_3901;
    end
    if (sel) begin
      lineBuffer_3903 <= lineBuffer_3902;
    end
    if (sel) begin
      lineBuffer_3904 <= lineBuffer_3903;
    end
    if (sel) begin
      lineBuffer_3905 <= lineBuffer_3904;
    end
    if (sel) begin
      lineBuffer_3906 <= lineBuffer_3905;
    end
    if (sel) begin
      lineBuffer_3907 <= lineBuffer_3906;
    end
    if (sel) begin
      lineBuffer_3908 <= lineBuffer_3907;
    end
    if (sel) begin
      lineBuffer_3909 <= lineBuffer_3908;
    end
    if (sel) begin
      lineBuffer_3910 <= lineBuffer_3909;
    end
    if (sel) begin
      lineBuffer_3911 <= lineBuffer_3910;
    end
    if (sel) begin
      lineBuffer_3912 <= lineBuffer_3911;
    end
    if (sel) begin
      lineBuffer_3913 <= lineBuffer_3912;
    end
    if (sel) begin
      lineBuffer_3914 <= lineBuffer_3913;
    end
    if (sel) begin
      lineBuffer_3915 <= lineBuffer_3914;
    end
    if (sel) begin
      lineBuffer_3916 <= lineBuffer_3915;
    end
    if (sel) begin
      lineBuffer_3917 <= lineBuffer_3916;
    end
    if (sel) begin
      lineBuffer_3918 <= lineBuffer_3917;
    end
    if (sel) begin
      lineBuffer_3919 <= lineBuffer_3918;
    end
    if (sel) begin
      lineBuffer_3920 <= lineBuffer_3919;
    end
    if (sel) begin
      lineBuffer_3921 <= lineBuffer_3920;
    end
    if (sel) begin
      lineBuffer_3922 <= lineBuffer_3921;
    end
    if (sel) begin
      lineBuffer_3923 <= lineBuffer_3922;
    end
    if (sel) begin
      lineBuffer_3924 <= lineBuffer_3923;
    end
    if (sel) begin
      lineBuffer_3925 <= lineBuffer_3924;
    end
    if (sel) begin
      lineBuffer_3926 <= lineBuffer_3925;
    end
    if (sel) begin
      lineBuffer_3927 <= lineBuffer_3926;
    end
    if (sel) begin
      lineBuffer_3928 <= lineBuffer_3927;
    end
    if (sel) begin
      lineBuffer_3929 <= lineBuffer_3928;
    end
    if (sel) begin
      lineBuffer_3930 <= lineBuffer_3929;
    end
    if (sel) begin
      lineBuffer_3931 <= lineBuffer_3930;
    end
    if (sel) begin
      lineBuffer_3932 <= lineBuffer_3931;
    end
    if (sel) begin
      lineBuffer_3933 <= lineBuffer_3932;
    end
    if (sel) begin
      lineBuffer_3934 <= lineBuffer_3933;
    end
    if (sel) begin
      lineBuffer_3935 <= lineBuffer_3934;
    end
    if (sel) begin
      lineBuffer_3936 <= lineBuffer_3935;
    end
    if (sel) begin
      lineBuffer_3937 <= lineBuffer_3936;
    end
    if (sel) begin
      lineBuffer_3938 <= lineBuffer_3937;
    end
    if (sel) begin
      lineBuffer_3939 <= lineBuffer_3938;
    end
    if (sel) begin
      lineBuffer_3940 <= lineBuffer_3939;
    end
    if (sel) begin
      lineBuffer_3941 <= lineBuffer_3940;
    end
    if (sel) begin
      lineBuffer_3942 <= lineBuffer_3941;
    end
    if (sel) begin
      lineBuffer_3943 <= lineBuffer_3942;
    end
    if (sel) begin
      lineBuffer_3944 <= lineBuffer_3943;
    end
    if (sel) begin
      lineBuffer_3945 <= lineBuffer_3944;
    end
    if (sel) begin
      lineBuffer_3946 <= lineBuffer_3945;
    end
    if (sel) begin
      lineBuffer_3947 <= lineBuffer_3946;
    end
    if (sel) begin
      lineBuffer_3948 <= lineBuffer_3947;
    end
    if (sel) begin
      lineBuffer_3949 <= lineBuffer_3948;
    end
    if (sel) begin
      lineBuffer_3950 <= lineBuffer_3949;
    end
    if (sel) begin
      lineBuffer_3951 <= lineBuffer_3950;
    end
    if (sel) begin
      lineBuffer_3952 <= lineBuffer_3951;
    end
    if (sel) begin
      lineBuffer_3953 <= lineBuffer_3952;
    end
    if (sel) begin
      lineBuffer_3954 <= lineBuffer_3953;
    end
    if (sel) begin
      lineBuffer_3955 <= lineBuffer_3954;
    end
    if (sel) begin
      lineBuffer_3956 <= lineBuffer_3955;
    end
    if (sel) begin
      lineBuffer_3957 <= lineBuffer_3956;
    end
    if (sel) begin
      lineBuffer_3958 <= lineBuffer_3957;
    end
    if (sel) begin
      lineBuffer_3959 <= lineBuffer_3958;
    end
    if (sel) begin
      lineBuffer_3960 <= lineBuffer_3959;
    end
    if (sel) begin
      lineBuffer_3961 <= lineBuffer_3960;
    end
    if (sel) begin
      lineBuffer_3962 <= lineBuffer_3961;
    end
    if (sel) begin
      lineBuffer_3963 <= lineBuffer_3962;
    end
    if (sel) begin
      lineBuffer_3964 <= lineBuffer_3963;
    end
    if (sel) begin
      lineBuffer_3965 <= lineBuffer_3964;
    end
    if (sel) begin
      lineBuffer_3966 <= lineBuffer_3965;
    end
    if (sel) begin
      lineBuffer_3967 <= lineBuffer_3966;
    end
    if (sel) begin
      lineBuffer_3968 <= lineBuffer_3967;
    end
    if (sel) begin
      lineBuffer_3969 <= lineBuffer_3968;
    end
    if (sel) begin
      lineBuffer_3970 <= lineBuffer_3969;
    end
    if (sel) begin
      lineBuffer_3971 <= lineBuffer_3970;
    end
    if (sel) begin
      lineBuffer_3972 <= lineBuffer_3971;
    end
    if (sel) begin
      lineBuffer_3973 <= lineBuffer_3972;
    end
    if (sel) begin
      lineBuffer_3974 <= lineBuffer_3973;
    end
    if (sel) begin
      lineBuffer_3975 <= lineBuffer_3974;
    end
    if (sel) begin
      lineBuffer_3976 <= lineBuffer_3975;
    end
    if (sel) begin
      lineBuffer_3977 <= lineBuffer_3976;
    end
    if (sel) begin
      lineBuffer_3978 <= lineBuffer_3977;
    end
    if (sel) begin
      lineBuffer_3979 <= lineBuffer_3978;
    end
    if (sel) begin
      lineBuffer_3980 <= lineBuffer_3979;
    end
    if (sel) begin
      lineBuffer_3981 <= lineBuffer_3980;
    end
    if (sel) begin
      lineBuffer_3982 <= lineBuffer_3981;
    end
    if (sel) begin
      lineBuffer_3983 <= lineBuffer_3982;
    end
    if (sel) begin
      lineBuffer_3984 <= lineBuffer_3983;
    end
    if (sel) begin
      lineBuffer_3985 <= lineBuffer_3984;
    end
    if (sel) begin
      lineBuffer_3986 <= lineBuffer_3985;
    end
    if (sel) begin
      lineBuffer_3987 <= lineBuffer_3986;
    end
    if (sel) begin
      lineBuffer_3988 <= lineBuffer_3987;
    end
    if (sel) begin
      lineBuffer_3989 <= lineBuffer_3988;
    end
    if (sel) begin
      lineBuffer_3990 <= lineBuffer_3989;
    end
    if (sel) begin
      lineBuffer_3991 <= lineBuffer_3990;
    end
    if (sel) begin
      lineBuffer_3992 <= lineBuffer_3991;
    end
    if (sel) begin
      lineBuffer_3993 <= lineBuffer_3992;
    end
    if (sel) begin
      lineBuffer_3994 <= lineBuffer_3993;
    end
    if (sel) begin
      lineBuffer_3995 <= lineBuffer_3994;
    end
    if (sel) begin
      lineBuffer_3996 <= lineBuffer_3995;
    end
    if (sel) begin
      lineBuffer_3997 <= lineBuffer_3996;
    end
    if (sel) begin
      lineBuffer_3998 <= lineBuffer_3997;
    end
    if (sel) begin
      lineBuffer_3999 <= lineBuffer_3998;
    end
    if (sel) begin
      lineBuffer_4000 <= lineBuffer_3999;
    end
    if (sel) begin
      lineBuffer_4001 <= lineBuffer_4000;
    end
    if (sel) begin
      lineBuffer_4002 <= lineBuffer_4001;
    end
    if (sel) begin
      lineBuffer_4003 <= lineBuffer_4002;
    end
    if (sel) begin
      lineBuffer_4004 <= lineBuffer_4003;
    end
    if (sel) begin
      lineBuffer_4005 <= lineBuffer_4004;
    end
    if (sel) begin
      lineBuffer_4006 <= lineBuffer_4005;
    end
    if (sel) begin
      lineBuffer_4007 <= lineBuffer_4006;
    end
    if (sel) begin
      lineBuffer_4008 <= lineBuffer_4007;
    end
    if (sel) begin
      lineBuffer_4009 <= lineBuffer_4008;
    end
    if (sel) begin
      lineBuffer_4010 <= lineBuffer_4009;
    end
    if (sel) begin
      lineBuffer_4011 <= lineBuffer_4010;
    end
    if (sel) begin
      lineBuffer_4012 <= lineBuffer_4011;
    end
    if (sel) begin
      lineBuffer_4013 <= lineBuffer_4012;
    end
    if (sel) begin
      lineBuffer_4014 <= lineBuffer_4013;
    end
    if (sel) begin
      lineBuffer_4015 <= lineBuffer_4014;
    end
    if (sel) begin
      lineBuffer_4016 <= lineBuffer_4015;
    end
    if (sel) begin
      lineBuffer_4017 <= lineBuffer_4016;
    end
    if (sel) begin
      lineBuffer_4018 <= lineBuffer_4017;
    end
    if (sel) begin
      lineBuffer_4019 <= lineBuffer_4018;
    end
    if (sel) begin
      lineBuffer_4020 <= lineBuffer_4019;
    end
    if (sel) begin
      lineBuffer_4021 <= lineBuffer_4020;
    end
    if (sel) begin
      lineBuffer_4022 <= lineBuffer_4021;
    end
    if (sel) begin
      lineBuffer_4023 <= lineBuffer_4022;
    end
    if (sel) begin
      lineBuffer_4024 <= lineBuffer_4023;
    end
    if (sel) begin
      lineBuffer_4025 <= lineBuffer_4024;
    end
    if (sel) begin
      lineBuffer_4026 <= lineBuffer_4025;
    end
    if (sel) begin
      lineBuffer_4027 <= lineBuffer_4026;
    end
    if (sel) begin
      lineBuffer_4028 <= lineBuffer_4027;
    end
    if (sel) begin
      lineBuffer_4029 <= lineBuffer_4028;
    end
    if (sel) begin
      lineBuffer_4030 <= lineBuffer_4029;
    end
    if (sel) begin
      lineBuffer_4031 <= lineBuffer_4030;
    end
    if (sel) begin
      lineBuffer_4032 <= lineBuffer_4031;
    end
    if (sel) begin
      lineBuffer_4033 <= lineBuffer_4032;
    end
    if (sel) begin
      lineBuffer_4034 <= lineBuffer_4033;
    end
    if (sel) begin
      lineBuffer_4035 <= lineBuffer_4034;
    end
    if (sel) begin
      lineBuffer_4036 <= lineBuffer_4035;
    end
    if (sel) begin
      lineBuffer_4037 <= lineBuffer_4036;
    end
    if (sel) begin
      lineBuffer_4038 <= lineBuffer_4037;
    end
    if (sel) begin
      lineBuffer_4039 <= lineBuffer_4038;
    end
    if (sel) begin
      lineBuffer_4040 <= lineBuffer_4039;
    end
    if (sel) begin
      lineBuffer_4041 <= lineBuffer_4040;
    end
    if (sel) begin
      lineBuffer_4042 <= lineBuffer_4041;
    end
    if (sel) begin
      lineBuffer_4043 <= lineBuffer_4042;
    end
    if (sel) begin
      lineBuffer_4044 <= lineBuffer_4043;
    end
    if (sel) begin
      lineBuffer_4045 <= lineBuffer_4044;
    end
    if (sel) begin
      lineBuffer_4046 <= lineBuffer_4045;
    end
    if (sel) begin
      lineBuffer_4047 <= lineBuffer_4046;
    end
    if (sel) begin
      lineBuffer_4048 <= lineBuffer_4047;
    end
    if (sel) begin
      lineBuffer_4049 <= lineBuffer_4048;
    end
    if (sel) begin
      lineBuffer_4050 <= lineBuffer_4049;
    end
    if (sel) begin
      lineBuffer_4051 <= lineBuffer_4050;
    end
    if (sel) begin
      lineBuffer_4052 <= lineBuffer_4051;
    end
    if (sel) begin
      lineBuffer_4053 <= lineBuffer_4052;
    end
    if (sel) begin
      lineBuffer_4054 <= lineBuffer_4053;
    end
    if (sel) begin
      lineBuffer_4055 <= lineBuffer_4054;
    end
    if (sel) begin
      lineBuffer_4056 <= lineBuffer_4055;
    end
    if (sel) begin
      lineBuffer_4057 <= lineBuffer_4056;
    end
    if (sel) begin
      lineBuffer_4058 <= lineBuffer_4057;
    end
    if (sel) begin
      lineBuffer_4059 <= lineBuffer_4058;
    end
    if (sel) begin
      lineBuffer_4060 <= lineBuffer_4059;
    end
    if (sel) begin
      lineBuffer_4061 <= lineBuffer_4060;
    end
    if (sel) begin
      lineBuffer_4062 <= lineBuffer_4061;
    end
    if (sel) begin
      lineBuffer_4063 <= lineBuffer_4062;
    end
    if (sel) begin
      lineBuffer_4064 <= lineBuffer_4063;
    end
    if (sel) begin
      lineBuffer_4065 <= lineBuffer_4064;
    end
    if (sel) begin
      lineBuffer_4066 <= lineBuffer_4065;
    end
    if (sel) begin
      lineBuffer_4067 <= lineBuffer_4066;
    end
    if (sel) begin
      lineBuffer_4068 <= lineBuffer_4067;
    end
    if (sel) begin
      lineBuffer_4069 <= lineBuffer_4068;
    end
    if (sel) begin
      lineBuffer_4070 <= lineBuffer_4069;
    end
    if (sel) begin
      lineBuffer_4071 <= lineBuffer_4070;
    end
    if (sel) begin
      lineBuffer_4072 <= lineBuffer_4071;
    end
    if (sel) begin
      lineBuffer_4073 <= lineBuffer_4072;
    end
    if (sel) begin
      lineBuffer_4074 <= lineBuffer_4073;
    end
    if (sel) begin
      lineBuffer_4075 <= lineBuffer_4074;
    end
    if (sel) begin
      lineBuffer_4076 <= lineBuffer_4075;
    end
    if (sel) begin
      lineBuffer_4077 <= lineBuffer_4076;
    end
    if (sel) begin
      lineBuffer_4078 <= lineBuffer_4077;
    end
    if (sel) begin
      lineBuffer_4079 <= lineBuffer_4078;
    end
    if (sel) begin
      lineBuffer_4080 <= lineBuffer_4079;
    end
    if (sel) begin
      lineBuffer_4081 <= lineBuffer_4080;
    end
    if (sel) begin
      lineBuffer_4082 <= lineBuffer_4081;
    end
    if (sel) begin
      lineBuffer_4083 <= lineBuffer_4082;
    end
    if (sel) begin
      lineBuffer_4084 <= lineBuffer_4083;
    end
    if (sel) begin
      lineBuffer_4085 <= lineBuffer_4084;
    end
    if (sel) begin
      lineBuffer_4086 <= lineBuffer_4085;
    end
    if (sel) begin
      lineBuffer_4087 <= lineBuffer_4086;
    end
    if (sel) begin
      lineBuffer_4088 <= lineBuffer_4087;
    end
    if (sel) begin
      lineBuffer_4089 <= lineBuffer_4088;
    end
    if (sel) begin
      lineBuffer_4090 <= lineBuffer_4089;
    end
    if (sel) begin
      lineBuffer_4091 <= lineBuffer_4090;
    end
    if (sel) begin
      lineBuffer_4092 <= lineBuffer_4091;
    end
    if (sel) begin
      lineBuffer_4093 <= lineBuffer_4092;
    end
    if (sel) begin
      lineBuffer_4094 <= lineBuffer_4093;
    end
    if (sel) begin
      lineBuffer_4095 <= lineBuffer_4094;
    end
    if (sel) begin
      lineBuffer_4096 <= lineBuffer_4095;
    end
    if (sel) begin
      lineBuffer_4097 <= lineBuffer_4096;
    end
    if (sel) begin
      lineBuffer_4098 <= lineBuffer_4097;
    end
    if (sel) begin
      lineBuffer_4099 <= lineBuffer_4098;
    end
    if (sel) begin
      lineBuffer_4100 <= lineBuffer_4099;
    end
    if (sel) begin
      lineBuffer_4101 <= lineBuffer_4100;
    end
    if (sel) begin
      lineBuffer_4102 <= lineBuffer_4101;
    end
    if (sel) begin
      lineBuffer_4103 <= lineBuffer_4102;
    end
    if (sel) begin
      lineBuffer_4104 <= lineBuffer_4103;
    end
    if (sel) begin
      lineBuffer_4105 <= lineBuffer_4104;
    end
    if (sel) begin
      lineBuffer_4106 <= lineBuffer_4105;
    end
    if (sel) begin
      lineBuffer_4107 <= lineBuffer_4106;
    end
    if (sel) begin
      lineBuffer_4108 <= lineBuffer_4107;
    end
    if (sel) begin
      lineBuffer_4109 <= lineBuffer_4108;
    end
    if (sel) begin
      lineBuffer_4110 <= lineBuffer_4109;
    end
    if (sel) begin
      lineBuffer_4111 <= lineBuffer_4110;
    end
    if (sel) begin
      lineBuffer_4112 <= lineBuffer_4111;
    end
    if (sel) begin
      lineBuffer_4113 <= lineBuffer_4112;
    end
    if (sel) begin
      lineBuffer_4114 <= lineBuffer_4113;
    end
    if (sel) begin
      lineBuffer_4115 <= lineBuffer_4114;
    end
    if (sel) begin
      lineBuffer_4116 <= lineBuffer_4115;
    end
    if (sel) begin
      lineBuffer_4117 <= lineBuffer_4116;
    end
    if (sel) begin
      lineBuffer_4118 <= lineBuffer_4117;
    end
    if (sel) begin
      lineBuffer_4119 <= lineBuffer_4118;
    end
    if (sel) begin
      lineBuffer_4120 <= lineBuffer_4119;
    end
    if (sel) begin
      lineBuffer_4121 <= lineBuffer_4120;
    end
    if (sel) begin
      lineBuffer_4122 <= lineBuffer_4121;
    end
    if (sel) begin
      lineBuffer_4123 <= lineBuffer_4122;
    end
    if (sel) begin
      lineBuffer_4124 <= lineBuffer_4123;
    end
    if (sel) begin
      lineBuffer_4125 <= lineBuffer_4124;
    end
    if (sel) begin
      lineBuffer_4126 <= lineBuffer_4125;
    end
    if (sel) begin
      lineBuffer_4127 <= lineBuffer_4126;
    end
    if (sel) begin
      lineBuffer_4128 <= lineBuffer_4127;
    end
    if (sel) begin
      lineBuffer_4129 <= lineBuffer_4128;
    end
    if (sel) begin
      lineBuffer_4130 <= lineBuffer_4129;
    end
    if (sel) begin
      lineBuffer_4131 <= lineBuffer_4130;
    end
    if (sel) begin
      lineBuffer_4132 <= lineBuffer_4131;
    end
    if (sel) begin
      lineBuffer_4133 <= lineBuffer_4132;
    end
    if (sel) begin
      lineBuffer_4134 <= lineBuffer_4133;
    end
    if (sel) begin
      lineBuffer_4135 <= lineBuffer_4134;
    end
    if (sel) begin
      lineBuffer_4136 <= lineBuffer_4135;
    end
    if (sel) begin
      lineBuffer_4137 <= lineBuffer_4136;
    end
    if (sel) begin
      lineBuffer_4138 <= lineBuffer_4137;
    end
    if (sel) begin
      lineBuffer_4139 <= lineBuffer_4138;
    end
    if (sel) begin
      lineBuffer_4140 <= lineBuffer_4139;
    end
    if (sel) begin
      lineBuffer_4141 <= lineBuffer_4140;
    end
    if (sel) begin
      lineBuffer_4142 <= lineBuffer_4141;
    end
    if (sel) begin
      lineBuffer_4143 <= lineBuffer_4142;
    end
    if (sel) begin
      lineBuffer_4144 <= lineBuffer_4143;
    end
    if (sel) begin
      lineBuffer_4145 <= lineBuffer_4144;
    end
    if (sel) begin
      lineBuffer_4146 <= lineBuffer_4145;
    end
    if (sel) begin
      lineBuffer_4147 <= lineBuffer_4146;
    end
    if (sel) begin
      lineBuffer_4148 <= lineBuffer_4147;
    end
    if (sel) begin
      lineBuffer_4149 <= lineBuffer_4148;
    end
    if (sel) begin
      lineBuffer_4150 <= lineBuffer_4149;
    end
    if (sel) begin
      lineBuffer_4151 <= lineBuffer_4150;
    end
    if (sel) begin
      lineBuffer_4152 <= lineBuffer_4151;
    end
    if (sel) begin
      lineBuffer_4153 <= lineBuffer_4152;
    end
    if (sel) begin
      lineBuffer_4154 <= lineBuffer_4153;
    end
    if (sel) begin
      lineBuffer_4155 <= lineBuffer_4154;
    end
    if (sel) begin
      lineBuffer_4156 <= lineBuffer_4155;
    end
    if (sel) begin
      lineBuffer_4157 <= lineBuffer_4156;
    end
    if (sel) begin
      lineBuffer_4158 <= lineBuffer_4157;
    end
    if (sel) begin
      lineBuffer_4159 <= lineBuffer_4158;
    end
    if (sel) begin
      lineBuffer_4160 <= lineBuffer_4159;
    end
    if (sel) begin
      lineBuffer_4161 <= lineBuffer_4160;
    end
    if (sel) begin
      lineBuffer_4162 <= lineBuffer_4161;
    end
    if (sel) begin
      lineBuffer_4163 <= lineBuffer_4162;
    end
    if (sel) begin
      lineBuffer_4164 <= lineBuffer_4163;
    end
    if (sel) begin
      lineBuffer_4165 <= lineBuffer_4164;
    end
    if (sel) begin
      lineBuffer_4166 <= lineBuffer_4165;
    end
    if (sel) begin
      lineBuffer_4167 <= lineBuffer_4166;
    end
    if (sel) begin
      lineBuffer_4168 <= lineBuffer_4167;
    end
    if (sel) begin
      lineBuffer_4169 <= lineBuffer_4168;
    end
    if (sel) begin
      lineBuffer_4170 <= lineBuffer_4169;
    end
    if (sel) begin
      lineBuffer_4171 <= lineBuffer_4170;
    end
    if (sel) begin
      lineBuffer_4172 <= lineBuffer_4171;
    end
    if (sel) begin
      lineBuffer_4173 <= lineBuffer_4172;
    end
    if (sel) begin
      lineBuffer_4174 <= lineBuffer_4173;
    end
    if (sel) begin
      lineBuffer_4175 <= lineBuffer_4174;
    end
    if (sel) begin
      lineBuffer_4176 <= lineBuffer_4175;
    end
    if (sel) begin
      lineBuffer_4177 <= lineBuffer_4176;
    end
    if (sel) begin
      lineBuffer_4178 <= lineBuffer_4177;
    end
    if (sel) begin
      lineBuffer_4179 <= lineBuffer_4178;
    end
    if (sel) begin
      lineBuffer_4180 <= lineBuffer_4179;
    end
    if (sel) begin
      lineBuffer_4181 <= lineBuffer_4180;
    end
    if (sel) begin
      lineBuffer_4182 <= lineBuffer_4181;
    end
    if (sel) begin
      lineBuffer_4183 <= lineBuffer_4182;
    end
    if (sel) begin
      lineBuffer_4184 <= lineBuffer_4183;
    end
    if (sel) begin
      lineBuffer_4185 <= lineBuffer_4184;
    end
    if (sel) begin
      lineBuffer_4186 <= lineBuffer_4185;
    end
    if (sel) begin
      lineBuffer_4187 <= lineBuffer_4186;
    end
    if (sel) begin
      lineBuffer_4188 <= lineBuffer_4187;
    end
    if (sel) begin
      lineBuffer_4189 <= lineBuffer_4188;
    end
    if (sel) begin
      lineBuffer_4190 <= lineBuffer_4189;
    end
    if (sel) begin
      lineBuffer_4191 <= lineBuffer_4190;
    end
    if (sel) begin
      lineBuffer_4192 <= lineBuffer_4191;
    end
    if (sel) begin
      lineBuffer_4193 <= lineBuffer_4192;
    end
    if (sel) begin
      lineBuffer_4194 <= lineBuffer_4193;
    end
    if (sel) begin
      lineBuffer_4195 <= lineBuffer_4194;
    end
    if (sel) begin
      lineBuffer_4196 <= lineBuffer_4195;
    end
    if (sel) begin
      lineBuffer_4197 <= lineBuffer_4196;
    end
    if (sel) begin
      lineBuffer_4198 <= lineBuffer_4197;
    end
    if (sel) begin
      lineBuffer_4199 <= lineBuffer_4198;
    end
    if (sel) begin
      lineBuffer_4200 <= lineBuffer_4199;
    end
    if (sel) begin
      lineBuffer_4201 <= lineBuffer_4200;
    end
    if (sel) begin
      lineBuffer_4202 <= lineBuffer_4201;
    end
    if (sel) begin
      lineBuffer_4203 <= lineBuffer_4202;
    end
    if (sel) begin
      lineBuffer_4204 <= lineBuffer_4203;
    end
    if (sel) begin
      lineBuffer_4205 <= lineBuffer_4204;
    end
    if (sel) begin
      lineBuffer_4206 <= lineBuffer_4205;
    end
    if (sel) begin
      lineBuffer_4207 <= lineBuffer_4206;
    end
    if (sel) begin
      lineBuffer_4208 <= lineBuffer_4207;
    end
    if (sel) begin
      lineBuffer_4209 <= lineBuffer_4208;
    end
    if (sel) begin
      lineBuffer_4210 <= lineBuffer_4209;
    end
    if (sel) begin
      lineBuffer_4211 <= lineBuffer_4210;
    end
    if (sel) begin
      lineBuffer_4212 <= lineBuffer_4211;
    end
    if (sel) begin
      lineBuffer_4213 <= lineBuffer_4212;
    end
    if (sel) begin
      lineBuffer_4214 <= lineBuffer_4213;
    end
    if (sel) begin
      lineBuffer_4215 <= lineBuffer_4214;
    end
    if (sel) begin
      lineBuffer_4216 <= lineBuffer_4215;
    end
    if (sel) begin
      lineBuffer_4217 <= lineBuffer_4216;
    end
    if (sel) begin
      lineBuffer_4218 <= lineBuffer_4217;
    end
    if (sel) begin
      lineBuffer_4219 <= lineBuffer_4218;
    end
    if (sel) begin
      lineBuffer_4220 <= lineBuffer_4219;
    end
    if (sel) begin
      lineBuffer_4221 <= lineBuffer_4220;
    end
    if (sel) begin
      lineBuffer_4222 <= lineBuffer_4221;
    end
    if (sel) begin
      lineBuffer_4223 <= lineBuffer_4222;
    end
    if (sel) begin
      lineBuffer_4224 <= lineBuffer_4223;
    end
    if (sel) begin
      lineBuffer_4225 <= lineBuffer_4224;
    end
    if (sel) begin
      lineBuffer_4226 <= lineBuffer_4225;
    end
    if (sel) begin
      lineBuffer_4227 <= lineBuffer_4226;
    end
    if (sel) begin
      lineBuffer_4228 <= lineBuffer_4227;
    end
    if (sel) begin
      lineBuffer_4229 <= lineBuffer_4228;
    end
    if (sel) begin
      lineBuffer_4230 <= lineBuffer_4229;
    end
    if (sel) begin
      lineBuffer_4231 <= lineBuffer_4230;
    end
    if (sel) begin
      lineBuffer_4232 <= lineBuffer_4231;
    end
    if (sel) begin
      lineBuffer_4233 <= lineBuffer_4232;
    end
    if (sel) begin
      lineBuffer_4234 <= lineBuffer_4233;
    end
    if (sel) begin
      lineBuffer_4235 <= lineBuffer_4234;
    end
    if (sel) begin
      lineBuffer_4236 <= lineBuffer_4235;
    end
    if (sel) begin
      lineBuffer_4237 <= lineBuffer_4236;
    end
    if (sel) begin
      lineBuffer_4238 <= lineBuffer_4237;
    end
    if (sel) begin
      lineBuffer_4239 <= lineBuffer_4238;
    end
    if (sel) begin
      lineBuffer_4240 <= lineBuffer_4239;
    end
    if (sel) begin
      lineBuffer_4241 <= lineBuffer_4240;
    end
    if (sel) begin
      lineBuffer_4242 <= lineBuffer_4241;
    end
    if (sel) begin
      lineBuffer_4243 <= lineBuffer_4242;
    end
    if (sel) begin
      lineBuffer_4244 <= lineBuffer_4243;
    end
    if (sel) begin
      lineBuffer_4245 <= lineBuffer_4244;
    end
    if (sel) begin
      lineBuffer_4246 <= lineBuffer_4245;
    end
    if (sel) begin
      lineBuffer_4247 <= lineBuffer_4246;
    end
    if (sel) begin
      lineBuffer_4248 <= lineBuffer_4247;
    end
    if (sel) begin
      lineBuffer_4249 <= lineBuffer_4248;
    end
    if (sel) begin
      lineBuffer_4250 <= lineBuffer_4249;
    end
    if (sel) begin
      lineBuffer_4251 <= lineBuffer_4250;
    end
    if (sel) begin
      lineBuffer_4252 <= lineBuffer_4251;
    end
    if (sel) begin
      lineBuffer_4253 <= lineBuffer_4252;
    end
    if (sel) begin
      lineBuffer_4254 <= lineBuffer_4253;
    end
    if (sel) begin
      lineBuffer_4255 <= lineBuffer_4254;
    end
    if (sel) begin
      lineBuffer_4256 <= lineBuffer_4255;
    end
    if (sel) begin
      lineBuffer_4257 <= lineBuffer_4256;
    end
    if (sel) begin
      lineBuffer_4258 <= lineBuffer_4257;
    end
    if (sel) begin
      lineBuffer_4259 <= lineBuffer_4258;
    end
    if (sel) begin
      lineBuffer_4260 <= lineBuffer_4259;
    end
    if (sel) begin
      lineBuffer_4261 <= lineBuffer_4260;
    end
    if (sel) begin
      lineBuffer_4262 <= lineBuffer_4261;
    end
    if (sel) begin
      lineBuffer_4263 <= lineBuffer_4262;
    end
    if (sel) begin
      lineBuffer_4264 <= lineBuffer_4263;
    end
    if (sel) begin
      lineBuffer_4265 <= lineBuffer_4264;
    end
    if (sel) begin
      lineBuffer_4266 <= lineBuffer_4265;
    end
    if (sel) begin
      lineBuffer_4267 <= lineBuffer_4266;
    end
    if (sel) begin
      lineBuffer_4268 <= lineBuffer_4267;
    end
    if (sel) begin
      lineBuffer_4269 <= lineBuffer_4268;
    end
    if (sel) begin
      lineBuffer_4270 <= lineBuffer_4269;
    end
    if (sel) begin
      lineBuffer_4271 <= lineBuffer_4270;
    end
    if (sel) begin
      lineBuffer_4272 <= lineBuffer_4271;
    end
    if (sel) begin
      lineBuffer_4273 <= lineBuffer_4272;
    end
    if (sel) begin
      lineBuffer_4274 <= lineBuffer_4273;
    end
    if (sel) begin
      lineBuffer_4275 <= lineBuffer_4274;
    end
    if (sel) begin
      lineBuffer_4276 <= lineBuffer_4275;
    end
    if (sel) begin
      lineBuffer_4277 <= lineBuffer_4276;
    end
    if (sel) begin
      lineBuffer_4278 <= lineBuffer_4277;
    end
    if (sel) begin
      lineBuffer_4279 <= lineBuffer_4278;
    end
    if (sel) begin
      lineBuffer_4280 <= lineBuffer_4279;
    end
    if (sel) begin
      lineBuffer_4281 <= lineBuffer_4280;
    end
    if (sel) begin
      lineBuffer_4282 <= lineBuffer_4281;
    end
    if (sel) begin
      lineBuffer_4283 <= lineBuffer_4282;
    end
    if (sel) begin
      lineBuffer_4284 <= lineBuffer_4283;
    end
    if (sel) begin
      lineBuffer_4285 <= lineBuffer_4284;
    end
    if (sel) begin
      lineBuffer_4286 <= lineBuffer_4285;
    end
    if (sel) begin
      lineBuffer_4287 <= lineBuffer_4286;
    end
    if (sel) begin
      lineBuffer_4288 <= lineBuffer_4287;
    end
    if (sel) begin
      lineBuffer_4289 <= lineBuffer_4288;
    end
    if (sel) begin
      lineBuffer_4290 <= lineBuffer_4289;
    end
    if (sel) begin
      lineBuffer_4291 <= lineBuffer_4290;
    end
    if (sel) begin
      lineBuffer_4292 <= lineBuffer_4291;
    end
    if (sel) begin
      lineBuffer_4293 <= lineBuffer_4292;
    end
    if (sel) begin
      lineBuffer_4294 <= lineBuffer_4293;
    end
    if (sel) begin
      lineBuffer_4295 <= lineBuffer_4294;
    end
    if (sel) begin
      lineBuffer_4296 <= lineBuffer_4295;
    end
    if (sel) begin
      lineBuffer_4297 <= lineBuffer_4296;
    end
    if (sel) begin
      lineBuffer_4298 <= lineBuffer_4297;
    end
    if (sel) begin
      lineBuffer_4299 <= lineBuffer_4298;
    end
    if (sel) begin
      lineBuffer_4300 <= lineBuffer_4299;
    end
    if (sel) begin
      lineBuffer_4301 <= lineBuffer_4300;
    end
    if (sel) begin
      lineBuffer_4302 <= lineBuffer_4301;
    end
    if (sel) begin
      lineBuffer_4303 <= lineBuffer_4302;
    end
    if (sel) begin
      lineBuffer_4304 <= lineBuffer_4303;
    end
    if (sel) begin
      lineBuffer_4305 <= lineBuffer_4304;
    end
    if (sel) begin
      lineBuffer_4306 <= lineBuffer_4305;
    end
    if (sel) begin
      lineBuffer_4307 <= lineBuffer_4306;
    end
    if (sel) begin
      lineBuffer_4308 <= lineBuffer_4307;
    end
    if (sel) begin
      lineBuffer_4309 <= lineBuffer_4308;
    end
    if (sel) begin
      lineBuffer_4310 <= lineBuffer_4309;
    end
    if (sel) begin
      lineBuffer_4311 <= lineBuffer_4310;
    end
    if (sel) begin
      lineBuffer_4312 <= lineBuffer_4311;
    end
    if (sel) begin
      lineBuffer_4313 <= lineBuffer_4312;
    end
    if (sel) begin
      lineBuffer_4314 <= lineBuffer_4313;
    end
    if (sel) begin
      lineBuffer_4315 <= lineBuffer_4314;
    end
    if (sel) begin
      lineBuffer_4316 <= lineBuffer_4315;
    end
    if (sel) begin
      lineBuffer_4317 <= lineBuffer_4316;
    end
    if (sel) begin
      lineBuffer_4318 <= lineBuffer_4317;
    end
    if (sel) begin
      lineBuffer_4319 <= lineBuffer_4318;
    end
    if (sel) begin
      lineBuffer_4320 <= lineBuffer_4319;
    end
    if (sel) begin
      lineBuffer_4321 <= lineBuffer_4320;
    end
    if (sel) begin
      lineBuffer_4322 <= lineBuffer_4321;
    end
    if (sel) begin
      lineBuffer_4323 <= lineBuffer_4322;
    end
    if (sel) begin
      lineBuffer_4324 <= lineBuffer_4323;
    end
    if (sel) begin
      lineBuffer_4325 <= lineBuffer_4324;
    end
    if (sel) begin
      lineBuffer_4326 <= lineBuffer_4325;
    end
    if (sel) begin
      lineBuffer_4327 <= lineBuffer_4326;
    end
    if (sel) begin
      lineBuffer_4328 <= lineBuffer_4327;
    end
    if (sel) begin
      lineBuffer_4329 <= lineBuffer_4328;
    end
    if (sel) begin
      lineBuffer_4330 <= lineBuffer_4329;
    end
    if (sel) begin
      lineBuffer_4331 <= lineBuffer_4330;
    end
    if (sel) begin
      lineBuffer_4332 <= lineBuffer_4331;
    end
    if (sel) begin
      lineBuffer_4333 <= lineBuffer_4332;
    end
    if (sel) begin
      lineBuffer_4334 <= lineBuffer_4333;
    end
    if (sel) begin
      lineBuffer_4335 <= lineBuffer_4334;
    end
    if (sel) begin
      lineBuffer_4336 <= lineBuffer_4335;
    end
    if (sel) begin
      lineBuffer_4337 <= lineBuffer_4336;
    end
    if (sel) begin
      lineBuffer_4338 <= lineBuffer_4337;
    end
    if (sel) begin
      lineBuffer_4339 <= lineBuffer_4338;
    end
    if (sel) begin
      lineBuffer_4340 <= lineBuffer_4339;
    end
    if (sel) begin
      lineBuffer_4341 <= lineBuffer_4340;
    end
    if (sel) begin
      lineBuffer_4342 <= lineBuffer_4341;
    end
    if (sel) begin
      lineBuffer_4343 <= lineBuffer_4342;
    end
    if (sel) begin
      lineBuffer_4344 <= lineBuffer_4343;
    end
    if (sel) begin
      lineBuffer_4345 <= lineBuffer_4344;
    end
    if (sel) begin
      lineBuffer_4346 <= lineBuffer_4345;
    end
    if (sel) begin
      lineBuffer_4347 <= lineBuffer_4346;
    end
    if (sel) begin
      lineBuffer_4348 <= lineBuffer_4347;
    end
    if (sel) begin
      lineBuffer_4349 <= lineBuffer_4348;
    end
    if (sel) begin
      lineBuffer_4350 <= lineBuffer_4349;
    end
    if (sel) begin
      lineBuffer_4351 <= lineBuffer_4350;
    end
    if (sel) begin
      lineBuffer_4352 <= lineBuffer_4351;
    end
    if (sel) begin
      lineBuffer_4353 <= lineBuffer_4352;
    end
    if (sel) begin
      lineBuffer_4354 <= lineBuffer_4353;
    end
    if (sel) begin
      lineBuffer_4355 <= lineBuffer_4354;
    end
    if (sel) begin
      lineBuffer_4356 <= lineBuffer_4355;
    end
    if (sel) begin
      lineBuffer_4357 <= lineBuffer_4356;
    end
    if (sel) begin
      lineBuffer_4358 <= lineBuffer_4357;
    end
    if (sel) begin
      lineBuffer_4359 <= lineBuffer_4358;
    end
    if (sel) begin
      lineBuffer_4360 <= lineBuffer_4359;
    end
    if (sel) begin
      lineBuffer_4361 <= lineBuffer_4360;
    end
    if (sel) begin
      lineBuffer_4362 <= lineBuffer_4361;
    end
    if (sel) begin
      lineBuffer_4363 <= lineBuffer_4362;
    end
    if (sel) begin
      lineBuffer_4364 <= lineBuffer_4363;
    end
    if (sel) begin
      lineBuffer_4365 <= lineBuffer_4364;
    end
    if (sel) begin
      lineBuffer_4366 <= lineBuffer_4365;
    end
    if (sel) begin
      lineBuffer_4367 <= lineBuffer_4366;
    end
    if (sel) begin
      lineBuffer_4368 <= lineBuffer_4367;
    end
    if (sel) begin
      lineBuffer_4369 <= lineBuffer_4368;
    end
    if (sel) begin
      lineBuffer_4370 <= lineBuffer_4369;
    end
    if (sel) begin
      lineBuffer_4371 <= lineBuffer_4370;
    end
    if (sel) begin
      lineBuffer_4372 <= lineBuffer_4371;
    end
    if (sel) begin
      lineBuffer_4373 <= lineBuffer_4372;
    end
    if (sel) begin
      lineBuffer_4374 <= lineBuffer_4373;
    end
    if (sel) begin
      lineBuffer_4375 <= lineBuffer_4374;
    end
    if (sel) begin
      lineBuffer_4376 <= lineBuffer_4375;
    end
    if (sel) begin
      lineBuffer_4377 <= lineBuffer_4376;
    end
    if (sel) begin
      lineBuffer_4378 <= lineBuffer_4377;
    end
    if (sel) begin
      lineBuffer_4379 <= lineBuffer_4378;
    end
    if (sel) begin
      lineBuffer_4380 <= lineBuffer_4379;
    end
    if (sel) begin
      lineBuffer_4381 <= lineBuffer_4380;
    end
    if (sel) begin
      lineBuffer_4382 <= lineBuffer_4381;
    end
    if (sel) begin
      lineBuffer_4383 <= lineBuffer_4382;
    end
    if (sel) begin
      lineBuffer_4384 <= lineBuffer_4383;
    end
    if (sel) begin
      lineBuffer_4385 <= lineBuffer_4384;
    end
    if (sel) begin
      lineBuffer_4386 <= lineBuffer_4385;
    end
    if (sel) begin
      lineBuffer_4387 <= lineBuffer_4386;
    end
    if (sel) begin
      lineBuffer_4388 <= lineBuffer_4387;
    end
    if (sel) begin
      lineBuffer_4389 <= lineBuffer_4388;
    end
    if (sel) begin
      lineBuffer_4390 <= lineBuffer_4389;
    end
    if (sel) begin
      lineBuffer_4391 <= lineBuffer_4390;
    end
    if (sel) begin
      lineBuffer_4392 <= lineBuffer_4391;
    end
    if (sel) begin
      lineBuffer_4393 <= lineBuffer_4392;
    end
    if (sel) begin
      lineBuffer_4394 <= lineBuffer_4393;
    end
    if (sel) begin
      lineBuffer_4395 <= lineBuffer_4394;
    end
    if (sel) begin
      lineBuffer_4396 <= lineBuffer_4395;
    end
    if (sel) begin
      lineBuffer_4397 <= lineBuffer_4396;
    end
    if (sel) begin
      lineBuffer_4398 <= lineBuffer_4397;
    end
    if (sel) begin
      lineBuffer_4399 <= lineBuffer_4398;
    end
    if (sel) begin
      lineBuffer_4400 <= lineBuffer_4399;
    end
    if (sel) begin
      lineBuffer_4401 <= lineBuffer_4400;
    end
    if (sel) begin
      lineBuffer_4402 <= lineBuffer_4401;
    end
    if (sel) begin
      lineBuffer_4403 <= lineBuffer_4402;
    end
    if (sel) begin
      lineBuffer_4404 <= lineBuffer_4403;
    end
    if (sel) begin
      lineBuffer_4405 <= lineBuffer_4404;
    end
    if (sel) begin
      lineBuffer_4406 <= lineBuffer_4405;
    end
    if (sel) begin
      lineBuffer_4407 <= lineBuffer_4406;
    end
    if (sel) begin
      lineBuffer_4408 <= lineBuffer_4407;
    end
    if (sel) begin
      lineBuffer_4409 <= lineBuffer_4408;
    end
    if (sel) begin
      lineBuffer_4410 <= lineBuffer_4409;
    end
    if (sel) begin
      lineBuffer_4411 <= lineBuffer_4410;
    end
    if (sel) begin
      lineBuffer_4412 <= lineBuffer_4411;
    end
    if (sel) begin
      lineBuffer_4413 <= lineBuffer_4412;
    end
    if (sel) begin
      lineBuffer_4414 <= lineBuffer_4413;
    end
    if (sel) begin
      lineBuffer_4415 <= lineBuffer_4414;
    end
    if (sel) begin
      lineBuffer_4416 <= lineBuffer_4415;
    end
    if (sel) begin
      lineBuffer_4417 <= lineBuffer_4416;
    end
    if (sel) begin
      lineBuffer_4418 <= lineBuffer_4417;
    end
    if (sel) begin
      lineBuffer_4419 <= lineBuffer_4418;
    end
    if (sel) begin
      lineBuffer_4420 <= lineBuffer_4419;
    end
    if (sel) begin
      lineBuffer_4421 <= lineBuffer_4420;
    end
    if (sel) begin
      lineBuffer_4422 <= lineBuffer_4421;
    end
    if (sel) begin
      lineBuffer_4423 <= lineBuffer_4422;
    end
    if (sel) begin
      lineBuffer_4424 <= lineBuffer_4423;
    end
    if (sel) begin
      lineBuffer_4425 <= lineBuffer_4424;
    end
    if (sel) begin
      lineBuffer_4426 <= lineBuffer_4425;
    end
    if (sel) begin
      lineBuffer_4427 <= lineBuffer_4426;
    end
    if (sel) begin
      lineBuffer_4428 <= lineBuffer_4427;
    end
    if (sel) begin
      lineBuffer_4429 <= lineBuffer_4428;
    end
    if (sel) begin
      lineBuffer_4430 <= lineBuffer_4429;
    end
    if (sel) begin
      lineBuffer_4431 <= lineBuffer_4430;
    end
    if (sel) begin
      lineBuffer_4432 <= lineBuffer_4431;
    end
    if (sel) begin
      lineBuffer_4433 <= lineBuffer_4432;
    end
    if (sel) begin
      lineBuffer_4434 <= lineBuffer_4433;
    end
    if (sel) begin
      lineBuffer_4435 <= lineBuffer_4434;
    end
    if (sel) begin
      lineBuffer_4436 <= lineBuffer_4435;
    end
    if (sel) begin
      lineBuffer_4437 <= lineBuffer_4436;
    end
    if (sel) begin
      lineBuffer_4438 <= lineBuffer_4437;
    end
    if (sel) begin
      lineBuffer_4439 <= lineBuffer_4438;
    end
    if (sel) begin
      lineBuffer_4440 <= lineBuffer_4439;
    end
    if (sel) begin
      lineBuffer_4441 <= lineBuffer_4440;
    end
    if (sel) begin
      lineBuffer_4442 <= lineBuffer_4441;
    end
    if (sel) begin
      lineBuffer_4443 <= lineBuffer_4442;
    end
    if (sel) begin
      lineBuffer_4444 <= lineBuffer_4443;
    end
    if (sel) begin
      lineBuffer_4445 <= lineBuffer_4444;
    end
    if (sel) begin
      lineBuffer_4446 <= lineBuffer_4445;
    end
    if (sel) begin
      lineBuffer_4447 <= lineBuffer_4446;
    end
    if (sel) begin
      lineBuffer_4448 <= lineBuffer_4447;
    end
    if (sel) begin
      lineBuffer_4449 <= lineBuffer_4448;
    end
    if (sel) begin
      lineBuffer_4450 <= lineBuffer_4449;
    end
    if (sel) begin
      lineBuffer_4451 <= lineBuffer_4450;
    end
    if (sel) begin
      lineBuffer_4452 <= lineBuffer_4451;
    end
    if (sel) begin
      lineBuffer_4453 <= lineBuffer_4452;
    end
    if (sel) begin
      lineBuffer_4454 <= lineBuffer_4453;
    end
    if (sel) begin
      lineBuffer_4455 <= lineBuffer_4454;
    end
    if (sel) begin
      lineBuffer_4456 <= lineBuffer_4455;
    end
    if (sel) begin
      lineBuffer_4457 <= lineBuffer_4456;
    end
    if (sel) begin
      lineBuffer_4458 <= lineBuffer_4457;
    end
    if (sel) begin
      lineBuffer_4459 <= lineBuffer_4458;
    end
    if (sel) begin
      lineBuffer_4460 <= lineBuffer_4459;
    end
    if (sel) begin
      lineBuffer_4461 <= lineBuffer_4460;
    end
    if (sel) begin
      lineBuffer_4462 <= lineBuffer_4461;
    end
    if (sel) begin
      lineBuffer_4463 <= lineBuffer_4462;
    end
    if (sel) begin
      lineBuffer_4464 <= lineBuffer_4463;
    end
    if (sel) begin
      lineBuffer_4465 <= lineBuffer_4464;
    end
    if (sel) begin
      lineBuffer_4466 <= lineBuffer_4465;
    end
    if (sel) begin
      lineBuffer_4467 <= lineBuffer_4466;
    end
    if (sel) begin
      lineBuffer_4468 <= lineBuffer_4467;
    end
    if (sel) begin
      lineBuffer_4469 <= lineBuffer_4468;
    end
    if (sel) begin
      lineBuffer_4470 <= lineBuffer_4469;
    end
    if (sel) begin
      lineBuffer_4471 <= lineBuffer_4470;
    end
    if (sel) begin
      lineBuffer_4472 <= lineBuffer_4471;
    end
    if (sel) begin
      lineBuffer_4473 <= lineBuffer_4472;
    end
    if (sel) begin
      lineBuffer_4474 <= lineBuffer_4473;
    end
    if (sel) begin
      lineBuffer_4475 <= lineBuffer_4474;
    end
    if (sel) begin
      lineBuffer_4476 <= lineBuffer_4475;
    end
    if (sel) begin
      lineBuffer_4477 <= lineBuffer_4476;
    end
    if (sel) begin
      lineBuffer_4478 <= lineBuffer_4477;
    end
    if (sel) begin
      lineBuffer_4479 <= lineBuffer_4478;
    end
    if (sel) begin
      lineBuffer_4480 <= lineBuffer_4479;
    end
    if (sel) begin
      lineBuffer_4481 <= lineBuffer_4480;
    end
    if (sel) begin
      lineBuffer_4482 <= lineBuffer_4481;
    end
    if (sel) begin
      lineBuffer_4483 <= lineBuffer_4482;
    end
    if (sel) begin
      lineBuffer_4484 <= lineBuffer_4483;
    end
    if (sel) begin
      lineBuffer_4485 <= lineBuffer_4484;
    end
    if (sel) begin
      lineBuffer_4486 <= lineBuffer_4485;
    end
    if (sel) begin
      lineBuffer_4487 <= lineBuffer_4486;
    end
    if (sel) begin
      lineBuffer_4488 <= lineBuffer_4487;
    end
    if (sel) begin
      lineBuffer_4489 <= lineBuffer_4488;
    end
    if (sel) begin
      lineBuffer_4490 <= lineBuffer_4489;
    end
    if (sel) begin
      lineBuffer_4491 <= lineBuffer_4490;
    end
    if (sel) begin
      lineBuffer_4492 <= lineBuffer_4491;
    end
    if (sel) begin
      lineBuffer_4493 <= lineBuffer_4492;
    end
    if (sel) begin
      lineBuffer_4494 <= lineBuffer_4493;
    end
    if (sel) begin
      lineBuffer_4495 <= lineBuffer_4494;
    end
    if (sel) begin
      lineBuffer_4496 <= lineBuffer_4495;
    end
    if (sel) begin
      lineBuffer_4497 <= lineBuffer_4496;
    end
    if (sel) begin
      lineBuffer_4498 <= lineBuffer_4497;
    end
    if (sel) begin
      lineBuffer_4499 <= lineBuffer_4498;
    end
    if (sel) begin
      lineBuffer_4500 <= lineBuffer_4499;
    end
    if (sel) begin
      lineBuffer_4501 <= lineBuffer_4500;
    end
    if (sel) begin
      lineBuffer_4502 <= lineBuffer_4501;
    end
    if (sel) begin
      lineBuffer_4503 <= lineBuffer_4502;
    end
    if (sel) begin
      lineBuffer_4504 <= lineBuffer_4503;
    end
    if (sel) begin
      lineBuffer_4505 <= lineBuffer_4504;
    end
    if (sel) begin
      lineBuffer_4506 <= lineBuffer_4505;
    end
    if (sel) begin
      lineBuffer_4507 <= lineBuffer_4506;
    end
    if (sel) begin
      lineBuffer_4508 <= lineBuffer_4507;
    end
    if (sel) begin
      lineBuffer_4509 <= lineBuffer_4508;
    end
    if (sel) begin
      lineBuffer_4510 <= lineBuffer_4509;
    end
    if (sel) begin
      lineBuffer_4511 <= lineBuffer_4510;
    end
    if (sel) begin
      lineBuffer_4512 <= lineBuffer_4511;
    end
    if (sel) begin
      lineBuffer_4513 <= lineBuffer_4512;
    end
    if (sel) begin
      lineBuffer_4514 <= lineBuffer_4513;
    end
    if (sel) begin
      lineBuffer_4515 <= lineBuffer_4514;
    end
    if (sel) begin
      lineBuffer_4516 <= lineBuffer_4515;
    end
    if (sel) begin
      lineBuffer_4517 <= lineBuffer_4516;
    end
    if (sel) begin
      lineBuffer_4518 <= lineBuffer_4517;
    end
    if (sel) begin
      lineBuffer_4519 <= lineBuffer_4518;
    end
    if (sel) begin
      lineBuffer_4520 <= lineBuffer_4519;
    end
    if (sel) begin
      lineBuffer_4521 <= lineBuffer_4520;
    end
    if (sel) begin
      lineBuffer_4522 <= lineBuffer_4521;
    end
    if (sel) begin
      lineBuffer_4523 <= lineBuffer_4522;
    end
    if (sel) begin
      lineBuffer_4524 <= lineBuffer_4523;
    end
    if (sel) begin
      lineBuffer_4525 <= lineBuffer_4524;
    end
    if (sel) begin
      lineBuffer_4526 <= lineBuffer_4525;
    end
    if (sel) begin
      lineBuffer_4527 <= lineBuffer_4526;
    end
    if (sel) begin
      lineBuffer_4528 <= lineBuffer_4527;
    end
    if (sel) begin
      lineBuffer_4529 <= lineBuffer_4528;
    end
    if (sel) begin
      lineBuffer_4530 <= lineBuffer_4529;
    end
    if (sel) begin
      lineBuffer_4531 <= lineBuffer_4530;
    end
    if (sel) begin
      lineBuffer_4532 <= lineBuffer_4531;
    end
    if (sel) begin
      lineBuffer_4533 <= lineBuffer_4532;
    end
    if (sel) begin
      lineBuffer_4534 <= lineBuffer_4533;
    end
    if (sel) begin
      lineBuffer_4535 <= lineBuffer_4534;
    end
    if (sel) begin
      lineBuffer_4536 <= lineBuffer_4535;
    end
    if (sel) begin
      lineBuffer_4537 <= lineBuffer_4536;
    end
    if (sel) begin
      lineBuffer_4538 <= lineBuffer_4537;
    end
    if (sel) begin
      lineBuffer_4539 <= lineBuffer_4538;
    end
    if (sel) begin
      lineBuffer_4540 <= lineBuffer_4539;
    end
    if (sel) begin
      lineBuffer_4541 <= lineBuffer_4540;
    end
    if (sel) begin
      lineBuffer_4542 <= lineBuffer_4541;
    end
    if (sel) begin
      lineBuffer_4543 <= lineBuffer_4542;
    end
    if (sel) begin
      lineBuffer_4544 <= lineBuffer_4543;
    end
    if (sel) begin
      lineBuffer_4545 <= lineBuffer_4544;
    end
    if (sel) begin
      lineBuffer_4546 <= lineBuffer_4545;
    end
    if (sel) begin
      lineBuffer_4547 <= lineBuffer_4546;
    end
    if (sel) begin
      lineBuffer_4548 <= lineBuffer_4547;
    end
    if (sel) begin
      lineBuffer_4549 <= lineBuffer_4548;
    end
    if (sel) begin
      lineBuffer_4550 <= lineBuffer_4549;
    end
    if (sel) begin
      lineBuffer_4551 <= lineBuffer_4550;
    end
    if (sel) begin
      lineBuffer_4552 <= lineBuffer_4551;
    end
    if (sel) begin
      lineBuffer_4553 <= lineBuffer_4552;
    end
    if (sel) begin
      lineBuffer_4554 <= lineBuffer_4553;
    end
    if (sel) begin
      lineBuffer_4555 <= lineBuffer_4554;
    end
    if (sel) begin
      lineBuffer_4556 <= lineBuffer_4555;
    end
    if (sel) begin
      lineBuffer_4557 <= lineBuffer_4556;
    end
    if (sel) begin
      lineBuffer_4558 <= lineBuffer_4557;
    end
    if (sel) begin
      lineBuffer_4559 <= lineBuffer_4558;
    end
    if (sel) begin
      lineBuffer_4560 <= lineBuffer_4559;
    end
    if (sel) begin
      lineBuffer_4561 <= lineBuffer_4560;
    end
    if (sel) begin
      lineBuffer_4562 <= lineBuffer_4561;
    end
    if (sel) begin
      lineBuffer_4563 <= lineBuffer_4562;
    end
    if (sel) begin
      lineBuffer_4564 <= lineBuffer_4563;
    end
    if (sel) begin
      lineBuffer_4565 <= lineBuffer_4564;
    end
    if (sel) begin
      lineBuffer_4566 <= lineBuffer_4565;
    end
    if (sel) begin
      lineBuffer_4567 <= lineBuffer_4566;
    end
    if (sel) begin
      lineBuffer_4568 <= lineBuffer_4567;
    end
    if (sel) begin
      lineBuffer_4569 <= lineBuffer_4568;
    end
    if (sel) begin
      lineBuffer_4570 <= lineBuffer_4569;
    end
    if (sel) begin
      lineBuffer_4571 <= lineBuffer_4570;
    end
    if (sel) begin
      lineBuffer_4572 <= lineBuffer_4571;
    end
    if (sel) begin
      lineBuffer_4573 <= lineBuffer_4572;
    end
    if (sel) begin
      lineBuffer_4574 <= lineBuffer_4573;
    end
    if (sel) begin
      lineBuffer_4575 <= lineBuffer_4574;
    end
    if (sel) begin
      lineBuffer_4576 <= lineBuffer_4575;
    end
    if (sel) begin
      lineBuffer_4577 <= lineBuffer_4576;
    end
    if (sel) begin
      lineBuffer_4578 <= lineBuffer_4577;
    end
    if (sel) begin
      lineBuffer_4579 <= lineBuffer_4578;
    end
    if (sel) begin
      lineBuffer_4580 <= lineBuffer_4579;
    end
    if (sel) begin
      lineBuffer_4581 <= lineBuffer_4580;
    end
    if (sel) begin
      lineBuffer_4582 <= lineBuffer_4581;
    end
    if (sel) begin
      lineBuffer_4583 <= lineBuffer_4582;
    end
    if (sel) begin
      lineBuffer_4584 <= lineBuffer_4583;
    end
    if (sel) begin
      lineBuffer_4585 <= lineBuffer_4584;
    end
    if (sel) begin
      lineBuffer_4586 <= lineBuffer_4585;
    end
    if (sel) begin
      lineBuffer_4587 <= lineBuffer_4586;
    end
    if (sel) begin
      lineBuffer_4588 <= lineBuffer_4587;
    end
    if (sel) begin
      lineBuffer_4589 <= lineBuffer_4588;
    end
    if (sel) begin
      lineBuffer_4590 <= lineBuffer_4589;
    end
    if (sel) begin
      lineBuffer_4591 <= lineBuffer_4590;
    end
    if (sel) begin
      lineBuffer_4592 <= lineBuffer_4591;
    end
    if (sel) begin
      lineBuffer_4593 <= lineBuffer_4592;
    end
    if (sel) begin
      lineBuffer_4594 <= lineBuffer_4593;
    end
    if (sel) begin
      lineBuffer_4595 <= lineBuffer_4594;
    end
    if (sel) begin
      lineBuffer_4596 <= lineBuffer_4595;
    end
    if (sel) begin
      lineBuffer_4597 <= lineBuffer_4596;
    end
    if (sel) begin
      lineBuffer_4598 <= lineBuffer_4597;
    end
    if (sel) begin
      lineBuffer_4599 <= lineBuffer_4598;
    end
    if (sel) begin
      lineBuffer_4600 <= lineBuffer_4599;
    end
    if (sel) begin
      lineBuffer_4601 <= lineBuffer_4600;
    end
    if (sel) begin
      lineBuffer_4602 <= lineBuffer_4601;
    end
    if (sel) begin
      lineBuffer_4603 <= lineBuffer_4602;
    end
    if (sel) begin
      lineBuffer_4604 <= lineBuffer_4603;
    end
    if (sel) begin
      lineBuffer_4605 <= lineBuffer_4604;
    end
    if (sel) begin
      lineBuffer_4606 <= lineBuffer_4605;
    end
    if (sel) begin
      lineBuffer_4607 <= lineBuffer_4606;
    end
    if (sel) begin
      lineBuffer_4608 <= lineBuffer_4607;
    end
    if (sel) begin
      lineBuffer_4609 <= lineBuffer_4608;
    end
    if (sel) begin
      lineBuffer_4610 <= lineBuffer_4609;
    end
    if (sel) begin
      lineBuffer_4611 <= lineBuffer_4610;
    end
    if (sel) begin
      lineBuffer_4612 <= lineBuffer_4611;
    end
    if (sel) begin
      lineBuffer_4613 <= lineBuffer_4612;
    end
    if (sel) begin
      lineBuffer_4614 <= lineBuffer_4613;
    end
    if (sel) begin
      lineBuffer_4615 <= lineBuffer_4614;
    end
    if (sel) begin
      lineBuffer_4616 <= lineBuffer_4615;
    end
    if (sel) begin
      lineBuffer_4617 <= lineBuffer_4616;
    end
    if (sel) begin
      lineBuffer_4618 <= lineBuffer_4617;
    end
    if (sel) begin
      lineBuffer_4619 <= lineBuffer_4618;
    end
    if (sel) begin
      lineBuffer_4620 <= lineBuffer_4619;
    end
    if (sel) begin
      lineBuffer_4621 <= lineBuffer_4620;
    end
    if (sel) begin
      lineBuffer_4622 <= lineBuffer_4621;
    end
    if (sel) begin
      lineBuffer_4623 <= lineBuffer_4622;
    end
    if (sel) begin
      lineBuffer_4624 <= lineBuffer_4623;
    end
    if (sel) begin
      lineBuffer_4625 <= lineBuffer_4624;
    end
    if (sel) begin
      lineBuffer_4626 <= lineBuffer_4625;
    end
    if (sel) begin
      lineBuffer_4627 <= lineBuffer_4626;
    end
    if (sel) begin
      lineBuffer_4628 <= lineBuffer_4627;
    end
    if (sel) begin
      lineBuffer_4629 <= lineBuffer_4628;
    end
    if (sel) begin
      lineBuffer_4630 <= lineBuffer_4629;
    end
    if (sel) begin
      lineBuffer_4631 <= lineBuffer_4630;
    end
    if (sel) begin
      lineBuffer_4632 <= lineBuffer_4631;
    end
    if (sel) begin
      lineBuffer_4633 <= lineBuffer_4632;
    end
    if (sel) begin
      lineBuffer_4634 <= lineBuffer_4633;
    end
    if (sel) begin
      lineBuffer_4635 <= lineBuffer_4634;
    end
    if (sel) begin
      lineBuffer_4636 <= lineBuffer_4635;
    end
    if (sel) begin
      lineBuffer_4637 <= lineBuffer_4636;
    end
    if (sel) begin
      lineBuffer_4638 <= lineBuffer_4637;
    end
    if (sel) begin
      lineBuffer_4639 <= lineBuffer_4638;
    end
    if (sel) begin
      lineBuffer_4640 <= lineBuffer_4639;
    end
    if (sel) begin
      lineBuffer_4641 <= lineBuffer_4640;
    end
    if (sel) begin
      lineBuffer_4642 <= lineBuffer_4641;
    end
    if (sel) begin
      lineBuffer_4643 <= lineBuffer_4642;
    end
    if (sel) begin
      lineBuffer_4644 <= lineBuffer_4643;
    end
    if (sel) begin
      lineBuffer_4645 <= lineBuffer_4644;
    end
    if (sel) begin
      lineBuffer_4646 <= lineBuffer_4645;
    end
    if (sel) begin
      lineBuffer_4647 <= lineBuffer_4646;
    end
    if (sel) begin
      lineBuffer_4648 <= lineBuffer_4647;
    end
    if (sel) begin
      lineBuffer_4649 <= lineBuffer_4648;
    end
    if (sel) begin
      lineBuffer_4650 <= lineBuffer_4649;
    end
    if (sel) begin
      lineBuffer_4651 <= lineBuffer_4650;
    end
    if (sel) begin
      lineBuffer_4652 <= lineBuffer_4651;
    end
    if (sel) begin
      lineBuffer_4653 <= lineBuffer_4652;
    end
    if (sel) begin
      lineBuffer_4654 <= lineBuffer_4653;
    end
    if (sel) begin
      lineBuffer_4655 <= lineBuffer_4654;
    end
    if (sel) begin
      lineBuffer_4656 <= lineBuffer_4655;
    end
    if (sel) begin
      lineBuffer_4657 <= lineBuffer_4656;
    end
    if (sel) begin
      lineBuffer_4658 <= lineBuffer_4657;
    end
    if (sel) begin
      lineBuffer_4659 <= lineBuffer_4658;
    end
    if (sel) begin
      lineBuffer_4660 <= lineBuffer_4659;
    end
    if (sel) begin
      lineBuffer_4661 <= lineBuffer_4660;
    end
    if (sel) begin
      lineBuffer_4662 <= lineBuffer_4661;
    end
    if (sel) begin
      lineBuffer_4663 <= lineBuffer_4662;
    end
    if (sel) begin
      lineBuffer_4664 <= lineBuffer_4663;
    end
    if (sel) begin
      lineBuffer_4665 <= lineBuffer_4664;
    end
    if (sel) begin
      lineBuffer_4666 <= lineBuffer_4665;
    end
    if (sel) begin
      lineBuffer_4667 <= lineBuffer_4666;
    end
    if (sel) begin
      lineBuffer_4668 <= lineBuffer_4667;
    end
    if (sel) begin
      lineBuffer_4669 <= lineBuffer_4668;
    end
    if (sel) begin
      lineBuffer_4670 <= lineBuffer_4669;
    end
    if (sel) begin
      lineBuffer_4671 <= lineBuffer_4670;
    end
    if (sel) begin
      lineBuffer_4672 <= lineBuffer_4671;
    end
    if (sel) begin
      lineBuffer_4673 <= lineBuffer_4672;
    end
    if (sel) begin
      lineBuffer_4674 <= lineBuffer_4673;
    end
    if (sel) begin
      lineBuffer_4675 <= lineBuffer_4674;
    end
    if (sel) begin
      lineBuffer_4676 <= lineBuffer_4675;
    end
    if (sel) begin
      lineBuffer_4677 <= lineBuffer_4676;
    end
    if (sel) begin
      lineBuffer_4678 <= lineBuffer_4677;
    end
    if (sel) begin
      lineBuffer_4679 <= lineBuffer_4678;
    end
    if (sel) begin
      lineBuffer_4680 <= lineBuffer_4679;
    end
    if (sel) begin
      lineBuffer_4681 <= lineBuffer_4680;
    end
    if (sel) begin
      lineBuffer_4682 <= lineBuffer_4681;
    end
    if (sel) begin
      lineBuffer_4683 <= lineBuffer_4682;
    end
    if (sel) begin
      lineBuffer_4684 <= lineBuffer_4683;
    end
    if (sel) begin
      lineBuffer_4685 <= lineBuffer_4684;
    end
    if (sel) begin
      lineBuffer_4686 <= lineBuffer_4685;
    end
    if (sel) begin
      lineBuffer_4687 <= lineBuffer_4686;
    end
    if (sel) begin
      lineBuffer_4688 <= lineBuffer_4687;
    end
    if (sel) begin
      lineBuffer_4689 <= lineBuffer_4688;
    end
    if (sel) begin
      lineBuffer_4690 <= lineBuffer_4689;
    end
    if (sel) begin
      lineBuffer_4691 <= lineBuffer_4690;
    end
    if (sel) begin
      lineBuffer_4692 <= lineBuffer_4691;
    end
    if (sel) begin
      lineBuffer_4693 <= lineBuffer_4692;
    end
    if (sel) begin
      lineBuffer_4694 <= lineBuffer_4693;
    end
    if (sel) begin
      lineBuffer_4695 <= lineBuffer_4694;
    end
    if (sel) begin
      lineBuffer_4696 <= lineBuffer_4695;
    end
    if (sel) begin
      lineBuffer_4697 <= lineBuffer_4696;
    end
    if (sel) begin
      lineBuffer_4698 <= lineBuffer_4697;
    end
    if (sel) begin
      lineBuffer_4699 <= lineBuffer_4698;
    end
    if (sel) begin
      lineBuffer_4700 <= lineBuffer_4699;
    end
    if (sel) begin
      lineBuffer_4701 <= lineBuffer_4700;
    end
    if (sel) begin
      lineBuffer_4702 <= lineBuffer_4701;
    end
    if (sel) begin
      lineBuffer_4703 <= lineBuffer_4702;
    end
    if (sel) begin
      lineBuffer_4704 <= lineBuffer_4703;
    end
    if (sel) begin
      lineBuffer_4705 <= lineBuffer_4704;
    end
    if (sel) begin
      lineBuffer_4706 <= lineBuffer_4705;
    end
    if (sel) begin
      lineBuffer_4707 <= lineBuffer_4706;
    end
    if (sel) begin
      lineBuffer_4708 <= lineBuffer_4707;
    end
    if (sel) begin
      lineBuffer_4709 <= lineBuffer_4708;
    end
    if (sel) begin
      lineBuffer_4710 <= lineBuffer_4709;
    end
    if (sel) begin
      lineBuffer_4711 <= lineBuffer_4710;
    end
    if (sel) begin
      lineBuffer_4712 <= lineBuffer_4711;
    end
    if (sel) begin
      lineBuffer_4713 <= lineBuffer_4712;
    end
    if (sel) begin
      lineBuffer_4714 <= lineBuffer_4713;
    end
    if (sel) begin
      lineBuffer_4715 <= lineBuffer_4714;
    end
    if (sel) begin
      lineBuffer_4716 <= lineBuffer_4715;
    end
    if (sel) begin
      lineBuffer_4717 <= lineBuffer_4716;
    end
    if (sel) begin
      lineBuffer_4718 <= lineBuffer_4717;
    end
    if (sel) begin
      lineBuffer_4719 <= lineBuffer_4718;
    end
    if (sel) begin
      lineBuffer_4720 <= lineBuffer_4719;
    end
    if (sel) begin
      lineBuffer_4721 <= lineBuffer_4720;
    end
    if (sel) begin
      lineBuffer_4722 <= lineBuffer_4721;
    end
    if (sel) begin
      lineBuffer_4723 <= lineBuffer_4722;
    end
    if (sel) begin
      lineBuffer_4724 <= lineBuffer_4723;
    end
    if (sel) begin
      lineBuffer_4725 <= lineBuffer_4724;
    end
    if (sel) begin
      lineBuffer_4726 <= lineBuffer_4725;
    end
    if (sel) begin
      lineBuffer_4727 <= lineBuffer_4726;
    end
    if (sel) begin
      lineBuffer_4728 <= lineBuffer_4727;
    end
    if (sel) begin
      lineBuffer_4729 <= lineBuffer_4728;
    end
    if (sel) begin
      lineBuffer_4730 <= lineBuffer_4729;
    end
    if (sel) begin
      lineBuffer_4731 <= lineBuffer_4730;
    end
    if (sel) begin
      lineBuffer_4732 <= lineBuffer_4731;
    end
    if (sel) begin
      lineBuffer_4733 <= lineBuffer_4732;
    end
    if (sel) begin
      lineBuffer_4734 <= lineBuffer_4733;
    end
    if (sel) begin
      lineBuffer_4735 <= lineBuffer_4734;
    end
    if (sel) begin
      lineBuffer_4736 <= lineBuffer_4735;
    end
    if (sel) begin
      lineBuffer_4737 <= lineBuffer_4736;
    end
    if (sel) begin
      lineBuffer_4738 <= lineBuffer_4737;
    end
    if (sel) begin
      lineBuffer_4739 <= lineBuffer_4738;
    end
    if (sel) begin
      lineBuffer_4740 <= lineBuffer_4739;
    end
    if (sel) begin
      lineBuffer_4741 <= lineBuffer_4740;
    end
    if (sel) begin
      lineBuffer_4742 <= lineBuffer_4741;
    end
    if (sel) begin
      lineBuffer_4743 <= lineBuffer_4742;
    end
    if (sel) begin
      lineBuffer_4744 <= lineBuffer_4743;
    end
    if (sel) begin
      lineBuffer_4745 <= lineBuffer_4744;
    end
    if (sel) begin
      lineBuffer_4746 <= lineBuffer_4745;
    end
    if (sel) begin
      lineBuffer_4747 <= lineBuffer_4746;
    end
    if (sel) begin
      lineBuffer_4748 <= lineBuffer_4747;
    end
    if (sel) begin
      lineBuffer_4749 <= lineBuffer_4748;
    end
    if (sel) begin
      lineBuffer_4750 <= lineBuffer_4749;
    end
    if (sel) begin
      lineBuffer_4751 <= lineBuffer_4750;
    end
    if (sel) begin
      lineBuffer_4752 <= lineBuffer_4751;
    end
    if (sel) begin
      lineBuffer_4753 <= lineBuffer_4752;
    end
    if (sel) begin
      lineBuffer_4754 <= lineBuffer_4753;
    end
    if (sel) begin
      lineBuffer_4755 <= lineBuffer_4754;
    end
    if (sel) begin
      lineBuffer_4756 <= lineBuffer_4755;
    end
    if (sel) begin
      lineBuffer_4757 <= lineBuffer_4756;
    end
    if (sel) begin
      lineBuffer_4758 <= lineBuffer_4757;
    end
    if (sel) begin
      lineBuffer_4759 <= lineBuffer_4758;
    end
    if (sel) begin
      lineBuffer_4760 <= lineBuffer_4759;
    end
    if (sel) begin
      lineBuffer_4761 <= lineBuffer_4760;
    end
    if (sel) begin
      lineBuffer_4762 <= lineBuffer_4761;
    end
    if (sel) begin
      lineBuffer_4763 <= lineBuffer_4762;
    end
    if (sel) begin
      lineBuffer_4764 <= lineBuffer_4763;
    end
    if (sel) begin
      lineBuffer_4765 <= lineBuffer_4764;
    end
    if (sel) begin
      lineBuffer_4766 <= lineBuffer_4765;
    end
    if (sel) begin
      lineBuffer_4767 <= lineBuffer_4766;
    end
    if (sel) begin
      lineBuffer_4768 <= lineBuffer_4767;
    end
    if (sel) begin
      lineBuffer_4769 <= lineBuffer_4768;
    end
    if (sel) begin
      lineBuffer_4770 <= lineBuffer_4769;
    end
    if (sel) begin
      lineBuffer_4771 <= lineBuffer_4770;
    end
    if (sel) begin
      lineBuffer_4772 <= lineBuffer_4771;
    end
    if (sel) begin
      lineBuffer_4773 <= lineBuffer_4772;
    end
    if (sel) begin
      lineBuffer_4774 <= lineBuffer_4773;
    end
    if (sel) begin
      lineBuffer_4775 <= lineBuffer_4774;
    end
    if (sel) begin
      lineBuffer_4776 <= lineBuffer_4775;
    end
    if (sel) begin
      lineBuffer_4777 <= lineBuffer_4776;
    end
    if (sel) begin
      lineBuffer_4778 <= lineBuffer_4777;
    end
    if (sel) begin
      lineBuffer_4779 <= lineBuffer_4778;
    end
    if (sel) begin
      lineBuffer_4780 <= lineBuffer_4779;
    end
    if (sel) begin
      lineBuffer_4781 <= lineBuffer_4780;
    end
    if (sel) begin
      lineBuffer_4782 <= lineBuffer_4781;
    end
    if (sel) begin
      lineBuffer_4783 <= lineBuffer_4782;
    end
    if (sel) begin
      lineBuffer_4784 <= lineBuffer_4783;
    end
    if (sel) begin
      lineBuffer_4785 <= lineBuffer_4784;
    end
    if (sel) begin
      lineBuffer_4786 <= lineBuffer_4785;
    end
    if (sel) begin
      lineBuffer_4787 <= lineBuffer_4786;
    end
    if (sel) begin
      lineBuffer_4788 <= lineBuffer_4787;
    end
    if (sel) begin
      lineBuffer_4789 <= lineBuffer_4788;
    end
    if (sel) begin
      lineBuffer_4790 <= lineBuffer_4789;
    end
    if (sel) begin
      lineBuffer_4791 <= lineBuffer_4790;
    end
    if (sel) begin
      lineBuffer_4792 <= lineBuffer_4791;
    end
    if (sel) begin
      lineBuffer_4793 <= lineBuffer_4792;
    end
    if (sel) begin
      lineBuffer_4794 <= lineBuffer_4793;
    end
    if (sel) begin
      lineBuffer_4795 <= lineBuffer_4794;
    end
    if (sel) begin
      lineBuffer_4796 <= lineBuffer_4795;
    end
    if (sel) begin
      lineBuffer_4797 <= lineBuffer_4796;
    end
    if (sel) begin
      lineBuffer_4798 <= lineBuffer_4797;
    end
    if (sel) begin
      lineBuffer_4799 <= lineBuffer_4798;
    end
    if (sel) begin
      lineBuffer_4800 <= lineBuffer_4799;
    end
    if (sel) begin
      lineBuffer_4801 <= lineBuffer_4800;
    end
    if (sel) begin
      lineBuffer_4802 <= lineBuffer_4801;
    end
    if (sel) begin
      lineBuffer_4803 <= lineBuffer_4802;
    end
    if (sel) begin
      lineBuffer_4804 <= lineBuffer_4803;
    end
    if (sel) begin
      lineBuffer_4805 <= lineBuffer_4804;
    end
    if (sel) begin
      lineBuffer_4806 <= lineBuffer_4805;
    end
    if (sel) begin
      lineBuffer_4807 <= lineBuffer_4806;
    end
    if (sel) begin
      lineBuffer_4808 <= lineBuffer_4807;
    end
    if (sel) begin
      lineBuffer_4809 <= lineBuffer_4808;
    end
    if (sel) begin
      lineBuffer_4810 <= lineBuffer_4809;
    end
    if (sel) begin
      lineBuffer_4811 <= lineBuffer_4810;
    end
    if (sel) begin
      lineBuffer_4812 <= lineBuffer_4811;
    end
    if (sel) begin
      lineBuffer_4813 <= lineBuffer_4812;
    end
    if (sel) begin
      lineBuffer_4814 <= lineBuffer_4813;
    end
    if (sel) begin
      lineBuffer_4815 <= lineBuffer_4814;
    end
    if (sel) begin
      lineBuffer_4816 <= lineBuffer_4815;
    end
    if (sel) begin
      lineBuffer_4817 <= lineBuffer_4816;
    end
    if (sel) begin
      lineBuffer_4818 <= lineBuffer_4817;
    end
    if (sel) begin
      lineBuffer_4819 <= lineBuffer_4818;
    end
    if (sel) begin
      lineBuffer_4820 <= lineBuffer_4819;
    end
    if (sel) begin
      lineBuffer_4821 <= lineBuffer_4820;
    end
    if (sel) begin
      lineBuffer_4822 <= lineBuffer_4821;
    end
    if (sel) begin
      lineBuffer_4823 <= lineBuffer_4822;
    end
    if (sel) begin
      lineBuffer_4824 <= lineBuffer_4823;
    end
    if (sel) begin
      lineBuffer_4825 <= lineBuffer_4824;
    end
    if (sel) begin
      lineBuffer_4826 <= lineBuffer_4825;
    end
    if (sel) begin
      lineBuffer_4827 <= lineBuffer_4826;
    end
    if (sel) begin
      lineBuffer_4828 <= lineBuffer_4827;
    end
    if (sel) begin
      lineBuffer_4829 <= lineBuffer_4828;
    end
    if (sel) begin
      lineBuffer_4830 <= lineBuffer_4829;
    end
    if (sel) begin
      lineBuffer_4831 <= lineBuffer_4830;
    end
    if (sel) begin
      lineBuffer_4832 <= lineBuffer_4831;
    end
    if (sel) begin
      lineBuffer_4833 <= lineBuffer_4832;
    end
    if (sel) begin
      lineBuffer_4834 <= lineBuffer_4833;
    end
    if (sel) begin
      lineBuffer_4835 <= lineBuffer_4834;
    end
    if (sel) begin
      lineBuffer_4836 <= lineBuffer_4835;
    end
    if (sel) begin
      lineBuffer_4837 <= lineBuffer_4836;
    end
    if (sel) begin
      lineBuffer_4838 <= lineBuffer_4837;
    end
    if (sel) begin
      lineBuffer_4839 <= lineBuffer_4838;
    end
    if (sel) begin
      lineBuffer_4840 <= lineBuffer_4839;
    end
    if (sel) begin
      lineBuffer_4841 <= lineBuffer_4840;
    end
    if (sel) begin
      lineBuffer_4842 <= lineBuffer_4841;
    end
    if (sel) begin
      lineBuffer_4843 <= lineBuffer_4842;
    end
    if (sel) begin
      lineBuffer_4844 <= lineBuffer_4843;
    end
    if (sel) begin
      lineBuffer_4845 <= lineBuffer_4844;
    end
    if (sel) begin
      lineBuffer_4846 <= lineBuffer_4845;
    end
    if (sel) begin
      lineBuffer_4847 <= lineBuffer_4846;
    end
    if (sel) begin
      lineBuffer_4848 <= lineBuffer_4847;
    end
    if (sel) begin
      lineBuffer_4849 <= lineBuffer_4848;
    end
    if (sel) begin
      lineBuffer_4850 <= lineBuffer_4849;
    end
    if (sel) begin
      lineBuffer_4851 <= lineBuffer_4850;
    end
    if (sel) begin
      lineBuffer_4852 <= lineBuffer_4851;
    end
    if (sel) begin
      lineBuffer_4853 <= lineBuffer_4852;
    end
    if (sel) begin
      lineBuffer_4854 <= lineBuffer_4853;
    end
    if (sel) begin
      lineBuffer_4855 <= lineBuffer_4854;
    end
    if (sel) begin
      lineBuffer_4856 <= lineBuffer_4855;
    end
    if (sel) begin
      lineBuffer_4857 <= lineBuffer_4856;
    end
    if (sel) begin
      lineBuffer_4858 <= lineBuffer_4857;
    end
    if (sel) begin
      lineBuffer_4859 <= lineBuffer_4858;
    end
    if (sel) begin
      lineBuffer_4860 <= lineBuffer_4859;
    end
    if (sel) begin
      lineBuffer_4861 <= lineBuffer_4860;
    end
    if (sel) begin
      lineBuffer_4862 <= lineBuffer_4861;
    end
    if (sel) begin
      lineBuffer_4863 <= lineBuffer_4862;
    end
    if (sel) begin
      lineBuffer_4864 <= lineBuffer_4863;
    end
    if (sel) begin
      lineBuffer_4865 <= lineBuffer_4864;
    end
    if (sel) begin
      lineBuffer_4866 <= lineBuffer_4865;
    end
    if (sel) begin
      lineBuffer_4867 <= lineBuffer_4866;
    end
    if (sel) begin
      lineBuffer_4868 <= lineBuffer_4867;
    end
    if (sel) begin
      lineBuffer_4869 <= lineBuffer_4868;
    end
    if (sel) begin
      lineBuffer_4870 <= lineBuffer_4869;
    end
    if (sel) begin
      lineBuffer_4871 <= lineBuffer_4870;
    end
    if (sel) begin
      lineBuffer_4872 <= lineBuffer_4871;
    end
    if (sel) begin
      lineBuffer_4873 <= lineBuffer_4872;
    end
    if (sel) begin
      lineBuffer_4874 <= lineBuffer_4873;
    end
    if (sel) begin
      lineBuffer_4875 <= lineBuffer_4874;
    end
    if (sel) begin
      lineBuffer_4876 <= lineBuffer_4875;
    end
    if (sel) begin
      lineBuffer_4877 <= lineBuffer_4876;
    end
    if (sel) begin
      lineBuffer_4878 <= lineBuffer_4877;
    end
    if (sel) begin
      lineBuffer_4879 <= lineBuffer_4878;
    end
    if (sel) begin
      lineBuffer_4880 <= lineBuffer_4879;
    end
    if (sel) begin
      lineBuffer_4881 <= lineBuffer_4880;
    end
    if (sel) begin
      lineBuffer_4882 <= lineBuffer_4881;
    end
    if (sel) begin
      lineBuffer_4883 <= lineBuffer_4882;
    end
    if (sel) begin
      lineBuffer_4884 <= lineBuffer_4883;
    end
    if (sel) begin
      lineBuffer_4885 <= lineBuffer_4884;
    end
    if (sel) begin
      lineBuffer_4886 <= lineBuffer_4885;
    end
    if (sel) begin
      lineBuffer_4887 <= lineBuffer_4886;
    end
    if (sel) begin
      lineBuffer_4888 <= lineBuffer_4887;
    end
    if (sel) begin
      lineBuffer_4889 <= lineBuffer_4888;
    end
    if (sel) begin
      lineBuffer_4890 <= lineBuffer_4889;
    end
    if (sel) begin
      lineBuffer_4891 <= lineBuffer_4890;
    end
    if (sel) begin
      lineBuffer_4892 <= lineBuffer_4891;
    end
    if (sel) begin
      lineBuffer_4893 <= lineBuffer_4892;
    end
    if (sel) begin
      lineBuffer_4894 <= lineBuffer_4893;
    end
    if (sel) begin
      lineBuffer_4895 <= lineBuffer_4894;
    end
    if (sel) begin
      lineBuffer_4896 <= lineBuffer_4895;
    end
    if (sel) begin
      lineBuffer_4897 <= lineBuffer_4896;
    end
    if (sel) begin
      lineBuffer_4898 <= lineBuffer_4897;
    end
    if (sel) begin
      lineBuffer_4899 <= lineBuffer_4898;
    end
    if (sel) begin
      lineBuffer_4900 <= lineBuffer_4899;
    end
    if (sel) begin
      lineBuffer_4901 <= lineBuffer_4900;
    end
    if (sel) begin
      lineBuffer_4902 <= lineBuffer_4901;
    end
    if (sel) begin
      lineBuffer_4903 <= lineBuffer_4902;
    end
    if (sel) begin
      lineBuffer_4904 <= lineBuffer_4903;
    end
    if (sel) begin
      lineBuffer_4905 <= lineBuffer_4904;
    end
    if (sel) begin
      lineBuffer_4906 <= lineBuffer_4905;
    end
    if (sel) begin
      lineBuffer_4907 <= lineBuffer_4906;
    end
    if (sel) begin
      lineBuffer_4908 <= lineBuffer_4907;
    end
    if (sel) begin
      lineBuffer_4909 <= lineBuffer_4908;
    end
    if (sel) begin
      lineBuffer_4910 <= lineBuffer_4909;
    end
    if (sel) begin
      lineBuffer_4911 <= lineBuffer_4910;
    end
    if (sel) begin
      lineBuffer_4912 <= lineBuffer_4911;
    end
    if (sel) begin
      lineBuffer_4913 <= lineBuffer_4912;
    end
    if (sel) begin
      lineBuffer_4914 <= lineBuffer_4913;
    end
    if (sel) begin
      lineBuffer_4915 <= lineBuffer_4914;
    end
    if (sel) begin
      lineBuffer_4916 <= lineBuffer_4915;
    end
    if (sel) begin
      lineBuffer_4917 <= lineBuffer_4916;
    end
    if (sel) begin
      lineBuffer_4918 <= lineBuffer_4917;
    end
    if (sel) begin
      lineBuffer_4919 <= lineBuffer_4918;
    end
    if (sel) begin
      lineBuffer_4920 <= lineBuffer_4919;
    end
    if (sel) begin
      lineBuffer_4921 <= lineBuffer_4920;
    end
    if (sel) begin
      lineBuffer_4922 <= lineBuffer_4921;
    end
    if (sel) begin
      lineBuffer_4923 <= lineBuffer_4922;
    end
    if (sel) begin
      lineBuffer_4924 <= lineBuffer_4923;
    end
    if (sel) begin
      lineBuffer_4925 <= lineBuffer_4924;
    end
    if (sel) begin
      lineBuffer_4926 <= lineBuffer_4925;
    end
    if (sel) begin
      lineBuffer_4927 <= lineBuffer_4926;
    end
    if (sel) begin
      lineBuffer_4928 <= lineBuffer_4927;
    end
    if (sel) begin
      lineBuffer_4929 <= lineBuffer_4928;
    end
    if (sel) begin
      lineBuffer_4930 <= lineBuffer_4929;
    end
    if (sel) begin
      lineBuffer_4931 <= lineBuffer_4930;
    end
    if (sel) begin
      lineBuffer_4932 <= lineBuffer_4931;
    end
    if (sel) begin
      lineBuffer_4933 <= lineBuffer_4932;
    end
    if (sel) begin
      lineBuffer_4934 <= lineBuffer_4933;
    end
    if (sel) begin
      lineBuffer_4935 <= lineBuffer_4934;
    end
    if (sel) begin
      lineBuffer_4936 <= lineBuffer_4935;
    end
    if (sel) begin
      lineBuffer_4937 <= lineBuffer_4936;
    end
    if (sel) begin
      lineBuffer_4938 <= lineBuffer_4937;
    end
    if (sel) begin
      lineBuffer_4939 <= lineBuffer_4938;
    end
    if (sel) begin
      lineBuffer_4940 <= lineBuffer_4939;
    end
    if (sel) begin
      lineBuffer_4941 <= lineBuffer_4940;
    end
    if (sel) begin
      lineBuffer_4942 <= lineBuffer_4941;
    end
    if (sel) begin
      lineBuffer_4943 <= lineBuffer_4942;
    end
    if (sel) begin
      lineBuffer_4944 <= lineBuffer_4943;
    end
    if (sel) begin
      lineBuffer_4945 <= lineBuffer_4944;
    end
    if (sel) begin
      lineBuffer_4946 <= lineBuffer_4945;
    end
    if (sel) begin
      lineBuffer_4947 <= lineBuffer_4946;
    end
    if (sel) begin
      lineBuffer_4948 <= lineBuffer_4947;
    end
    if (sel) begin
      lineBuffer_4949 <= lineBuffer_4948;
    end
    if (sel) begin
      lineBuffer_4950 <= lineBuffer_4949;
    end
    if (sel) begin
      lineBuffer_4951 <= lineBuffer_4950;
    end
    if (sel) begin
      lineBuffer_4952 <= lineBuffer_4951;
    end
    if (sel) begin
      lineBuffer_4953 <= lineBuffer_4952;
    end
    if (sel) begin
      lineBuffer_4954 <= lineBuffer_4953;
    end
    if (sel) begin
      lineBuffer_4955 <= lineBuffer_4954;
    end
    if (sel) begin
      lineBuffer_4956 <= lineBuffer_4955;
    end
    if (sel) begin
      lineBuffer_4957 <= lineBuffer_4956;
    end
    if (sel) begin
      lineBuffer_4958 <= lineBuffer_4957;
    end
    if (sel) begin
      lineBuffer_4959 <= lineBuffer_4958;
    end
    if (sel) begin
      lineBuffer_4960 <= lineBuffer_4959;
    end
    if (sel) begin
      lineBuffer_4961 <= lineBuffer_4960;
    end
    if (sel) begin
      lineBuffer_4962 <= lineBuffer_4961;
    end
    if (sel) begin
      lineBuffer_4963 <= lineBuffer_4962;
    end
    if (sel) begin
      lineBuffer_4964 <= lineBuffer_4963;
    end
    if (sel) begin
      lineBuffer_4965 <= lineBuffer_4964;
    end
    if (sel) begin
      lineBuffer_4966 <= lineBuffer_4965;
    end
    if (sel) begin
      lineBuffer_4967 <= lineBuffer_4966;
    end
    if (sel) begin
      lineBuffer_4968 <= lineBuffer_4967;
    end
    if (sel) begin
      lineBuffer_4969 <= lineBuffer_4968;
    end
    if (sel) begin
      lineBuffer_4970 <= lineBuffer_4969;
    end
    if (sel) begin
      lineBuffer_4971 <= lineBuffer_4970;
    end
    if (sel) begin
      lineBuffer_4972 <= lineBuffer_4971;
    end
    if (sel) begin
      lineBuffer_4973 <= lineBuffer_4972;
    end
    if (sel) begin
      lineBuffer_4974 <= lineBuffer_4973;
    end
    if (sel) begin
      lineBuffer_4975 <= lineBuffer_4974;
    end
    if (sel) begin
      lineBuffer_4976 <= lineBuffer_4975;
    end
    if (sel) begin
      lineBuffer_4977 <= lineBuffer_4976;
    end
    if (sel) begin
      lineBuffer_4978 <= lineBuffer_4977;
    end
    if (sel) begin
      lineBuffer_4979 <= lineBuffer_4978;
    end
    if (sel) begin
      lineBuffer_4980 <= lineBuffer_4979;
    end
    if (sel) begin
      lineBuffer_4981 <= lineBuffer_4980;
    end
    if (sel) begin
      lineBuffer_4982 <= lineBuffer_4981;
    end
    if (sel) begin
      lineBuffer_4983 <= lineBuffer_4982;
    end
    if (sel) begin
      lineBuffer_4984 <= lineBuffer_4983;
    end
    if (sel) begin
      lineBuffer_4985 <= lineBuffer_4984;
    end
    if (sel) begin
      lineBuffer_4986 <= lineBuffer_4985;
    end
    if (sel) begin
      lineBuffer_4987 <= lineBuffer_4986;
    end
    if (sel) begin
      lineBuffer_4988 <= lineBuffer_4987;
    end
    if (sel) begin
      lineBuffer_4989 <= lineBuffer_4988;
    end
    if (sel) begin
      lineBuffer_4990 <= lineBuffer_4989;
    end
    if (sel) begin
      lineBuffer_4991 <= lineBuffer_4990;
    end
    if (sel) begin
      lineBuffer_4992 <= lineBuffer_4991;
    end
    if (sel) begin
      lineBuffer_4993 <= lineBuffer_4992;
    end
    if (sel) begin
      lineBuffer_4994 <= lineBuffer_4993;
    end
    if (sel) begin
      lineBuffer_4995 <= lineBuffer_4994;
    end
    if (sel) begin
      lineBuffer_4996 <= lineBuffer_4995;
    end
    if (sel) begin
      lineBuffer_4997 <= lineBuffer_4996;
    end
    if (sel) begin
      lineBuffer_4998 <= lineBuffer_4997;
    end
    if (sel) begin
      lineBuffer_4999 <= lineBuffer_4998;
    end
    if (sel) begin
      lineBuffer_5000 <= lineBuffer_4999;
    end
    if (sel) begin
      lineBuffer_5001 <= lineBuffer_5000;
    end
    if (sel) begin
      lineBuffer_5002 <= lineBuffer_5001;
    end
    if (sel) begin
      lineBuffer_5003 <= lineBuffer_5002;
    end
    if (sel) begin
      lineBuffer_5004 <= lineBuffer_5003;
    end
    if (sel) begin
      lineBuffer_5005 <= lineBuffer_5004;
    end
    if (sel) begin
      lineBuffer_5006 <= lineBuffer_5005;
    end
    if (sel) begin
      lineBuffer_5007 <= lineBuffer_5006;
    end
    if (sel) begin
      lineBuffer_5008 <= lineBuffer_5007;
    end
    if (sel) begin
      lineBuffer_5009 <= lineBuffer_5008;
    end
    if (sel) begin
      lineBuffer_5010 <= lineBuffer_5009;
    end
    if (sel) begin
      lineBuffer_5011 <= lineBuffer_5010;
    end
    if (sel) begin
      lineBuffer_5012 <= lineBuffer_5011;
    end
    if (sel) begin
      lineBuffer_5013 <= lineBuffer_5012;
    end
    if (sel) begin
      lineBuffer_5014 <= lineBuffer_5013;
    end
    if (sel) begin
      lineBuffer_5015 <= lineBuffer_5014;
    end
    if (sel) begin
      lineBuffer_5016 <= lineBuffer_5015;
    end
    if (sel) begin
      lineBuffer_5017 <= lineBuffer_5016;
    end
    if (sel) begin
      lineBuffer_5018 <= lineBuffer_5017;
    end
    if (sel) begin
      lineBuffer_5019 <= lineBuffer_5018;
    end
    if (sel) begin
      lineBuffer_5020 <= lineBuffer_5019;
    end
    if (sel) begin
      lineBuffer_5021 <= lineBuffer_5020;
    end
    if (sel) begin
      lineBuffer_5022 <= lineBuffer_5021;
    end
    if (sel) begin
      lineBuffer_5023 <= lineBuffer_5022;
    end
    if (sel) begin
      lineBuffer_5024 <= lineBuffer_5023;
    end
    if (sel) begin
      lineBuffer_5025 <= lineBuffer_5024;
    end
    if (sel) begin
      lineBuffer_5026 <= lineBuffer_5025;
    end
    if (sel) begin
      lineBuffer_5027 <= lineBuffer_5026;
    end
    if (sel) begin
      lineBuffer_5028 <= lineBuffer_5027;
    end
    if (sel) begin
      lineBuffer_5029 <= lineBuffer_5028;
    end
    if (sel) begin
      lineBuffer_5030 <= lineBuffer_5029;
    end
    if (sel) begin
      lineBuffer_5031 <= lineBuffer_5030;
    end
    if (sel) begin
      lineBuffer_5032 <= lineBuffer_5031;
    end
    if (sel) begin
      lineBuffer_5033 <= lineBuffer_5032;
    end
    if (sel) begin
      lineBuffer_5034 <= lineBuffer_5033;
    end
    if (sel) begin
      lineBuffer_5035 <= lineBuffer_5034;
    end
    if (sel) begin
      lineBuffer_5036 <= lineBuffer_5035;
    end
    if (sel) begin
      lineBuffer_5037 <= lineBuffer_5036;
    end
    if (sel) begin
      lineBuffer_5038 <= lineBuffer_5037;
    end
    if (sel) begin
      lineBuffer_5039 <= lineBuffer_5038;
    end
    if (sel) begin
      lineBuffer_5040 <= lineBuffer_5039;
    end
    if (sel) begin
      lineBuffer_5041 <= lineBuffer_5040;
    end
    if (sel) begin
      lineBuffer_5042 <= lineBuffer_5041;
    end
    if (sel) begin
      lineBuffer_5043 <= lineBuffer_5042;
    end
    if (sel) begin
      lineBuffer_5044 <= lineBuffer_5043;
    end
    if (sel) begin
      lineBuffer_5045 <= lineBuffer_5044;
    end
    if (sel) begin
      lineBuffer_5046 <= lineBuffer_5045;
    end
    if (sel) begin
      lineBuffer_5047 <= lineBuffer_5046;
    end
    if (sel) begin
      lineBuffer_5048 <= lineBuffer_5047;
    end
    if (sel) begin
      lineBuffer_5049 <= lineBuffer_5048;
    end
    if (sel) begin
      lineBuffer_5050 <= lineBuffer_5049;
    end
    if (sel) begin
      lineBuffer_5051 <= lineBuffer_5050;
    end
    if (sel) begin
      lineBuffer_5052 <= lineBuffer_5051;
    end
    if (sel) begin
      lineBuffer_5053 <= lineBuffer_5052;
    end
    if (sel) begin
      lineBuffer_5054 <= lineBuffer_5053;
    end
    if (sel) begin
      lineBuffer_5055 <= lineBuffer_5054;
    end
    if (sel) begin
      lineBuffer_5056 <= lineBuffer_5055;
    end
    if (sel) begin
      lineBuffer_5057 <= lineBuffer_5056;
    end
    if (sel) begin
      lineBuffer_5058 <= lineBuffer_5057;
    end
    if (sel) begin
      lineBuffer_5059 <= lineBuffer_5058;
    end
    if (sel) begin
      lineBuffer_5060 <= lineBuffer_5059;
    end
    if (sel) begin
      lineBuffer_5061 <= lineBuffer_5060;
    end
    if (sel) begin
      lineBuffer_5062 <= lineBuffer_5061;
    end
    if (sel) begin
      lineBuffer_5063 <= lineBuffer_5062;
    end
    if (sel) begin
      lineBuffer_5064 <= lineBuffer_5063;
    end
    if (sel) begin
      lineBuffer_5065 <= lineBuffer_5064;
    end
    if (sel) begin
      lineBuffer_5066 <= lineBuffer_5065;
    end
    if (sel) begin
      lineBuffer_5067 <= lineBuffer_5066;
    end
    if (sel) begin
      lineBuffer_5068 <= lineBuffer_5067;
    end
    if (sel) begin
      lineBuffer_5069 <= lineBuffer_5068;
    end
    if (sel) begin
      lineBuffer_5070 <= lineBuffer_5069;
    end
    if (sel) begin
      lineBuffer_5071 <= lineBuffer_5070;
    end
    if (sel) begin
      lineBuffer_5072 <= lineBuffer_5071;
    end
    if (sel) begin
      lineBuffer_5073 <= lineBuffer_5072;
    end
    if (sel) begin
      lineBuffer_5074 <= lineBuffer_5073;
    end
    if (sel) begin
      lineBuffer_5075 <= lineBuffer_5074;
    end
    if (sel) begin
      lineBuffer_5076 <= lineBuffer_5075;
    end
    if (sel) begin
      lineBuffer_5077 <= lineBuffer_5076;
    end
    if (sel) begin
      lineBuffer_5078 <= lineBuffer_5077;
    end
    if (sel) begin
      lineBuffer_5079 <= lineBuffer_5078;
    end
    if (sel) begin
      lineBuffer_5080 <= lineBuffer_5079;
    end
    if (sel) begin
      lineBuffer_5081 <= lineBuffer_5080;
    end
    if (sel) begin
      lineBuffer_5082 <= lineBuffer_5081;
    end
    if (sel) begin
      lineBuffer_5083 <= lineBuffer_5082;
    end
    if (sel) begin
      lineBuffer_5084 <= lineBuffer_5083;
    end
    if (sel) begin
      lineBuffer_5085 <= lineBuffer_5084;
    end
    if (sel) begin
      lineBuffer_5086 <= lineBuffer_5085;
    end
    if (sel) begin
      lineBuffer_5087 <= lineBuffer_5086;
    end
    if (sel) begin
      lineBuffer_5088 <= lineBuffer_5087;
    end
    if (sel) begin
      lineBuffer_5089 <= lineBuffer_5088;
    end
    if (sel) begin
      lineBuffer_5090 <= lineBuffer_5089;
    end
    if (sel) begin
      lineBuffer_5091 <= lineBuffer_5090;
    end
    if (sel) begin
      lineBuffer_5092 <= lineBuffer_5091;
    end
    if (sel) begin
      lineBuffer_5093 <= lineBuffer_5092;
    end
    if (sel) begin
      lineBuffer_5094 <= lineBuffer_5093;
    end
    if (sel) begin
      lineBuffer_5095 <= lineBuffer_5094;
    end
    if (sel) begin
      lineBuffer_5096 <= lineBuffer_5095;
    end
    if (sel) begin
      lineBuffer_5097 <= lineBuffer_5096;
    end
    if (sel) begin
      lineBuffer_5098 <= lineBuffer_5097;
    end
    if (sel) begin
      lineBuffer_5099 <= lineBuffer_5098;
    end
    if (sel) begin
      lineBuffer_5100 <= lineBuffer_5099;
    end
    if (sel) begin
      lineBuffer_5101 <= lineBuffer_5100;
    end
    if (sel) begin
      lineBuffer_5102 <= lineBuffer_5101;
    end
    if (sel) begin
      lineBuffer_5103 <= lineBuffer_5102;
    end
    if (sel) begin
      lineBuffer_5104 <= lineBuffer_5103;
    end
    if (sel) begin
      lineBuffer_5105 <= lineBuffer_5104;
    end
    if (sel) begin
      lineBuffer_5106 <= lineBuffer_5105;
    end
    if (sel) begin
      lineBuffer_5107 <= lineBuffer_5106;
    end
    if (sel) begin
      lineBuffer_5108 <= lineBuffer_5107;
    end
    if (sel) begin
      lineBuffer_5109 <= lineBuffer_5108;
    end
    if (sel) begin
      lineBuffer_5110 <= lineBuffer_5109;
    end
    if (sel) begin
      lineBuffer_5111 <= lineBuffer_5110;
    end
    if (sel) begin
      lineBuffer_5112 <= lineBuffer_5111;
    end
    if (sel) begin
      lineBuffer_5113 <= lineBuffer_5112;
    end
    if (sel) begin
      lineBuffer_5114 <= lineBuffer_5113;
    end
    if (sel) begin
      lineBuffer_5115 <= lineBuffer_5114;
    end
    if (sel) begin
      lineBuffer_5116 <= lineBuffer_5115;
    end
    if (sel) begin
      lineBuffer_5117 <= lineBuffer_5116;
    end
    if (sel) begin
      lineBuffer_5118 <= lineBuffer_5117;
    end
    if (sel) begin
      lineBuffer_5119 <= lineBuffer_5118;
    end
    if (sel) begin
      lineBuffer_5120 <= lineBuffer_5119;
    end
    if (sel) begin
      lineBuffer_5121 <= lineBuffer_5120;
    end
    if (sel) begin
      lineBuffer_5122 <= lineBuffer_5121;
    end
    if (sel) begin
      lineBuffer_5123 <= lineBuffer_5122;
    end
    if (sel) begin
      lineBuffer_5124 <= lineBuffer_5123;
    end
    if (sel) begin
      lineBuffer_5125 <= lineBuffer_5124;
    end
    if (sel) begin
      lineBuffer_5126 <= lineBuffer_5125;
    end
    if (sel) begin
      lineBuffer_5127 <= lineBuffer_5126;
    end
    if (sel) begin
      lineBuffer_5128 <= lineBuffer_5127;
    end
    if (sel) begin
      lineBuffer_5129 <= lineBuffer_5128;
    end
    if (sel) begin
      lineBuffer_5130 <= lineBuffer_5129;
    end
    if (sel) begin
      lineBuffer_5131 <= lineBuffer_5130;
    end
    if (sel) begin
      lineBuffer_5132 <= lineBuffer_5131;
    end
    if (sel) begin
      lineBuffer_5133 <= lineBuffer_5132;
    end
    if (sel) begin
      lineBuffer_5134 <= lineBuffer_5133;
    end
    if (sel) begin
      lineBuffer_5135 <= lineBuffer_5134;
    end
    if (sel) begin
      lineBuffer_5136 <= lineBuffer_5135;
    end
    if (sel) begin
      lineBuffer_5137 <= lineBuffer_5136;
    end
    if (sel) begin
      lineBuffer_5138 <= lineBuffer_5137;
    end
    if (sel) begin
      lineBuffer_5139 <= lineBuffer_5138;
    end
    if (sel) begin
      lineBuffer_5140 <= lineBuffer_5139;
    end
    if (sel) begin
      lineBuffer_5141 <= lineBuffer_5140;
    end
    if (sel) begin
      lineBuffer_5142 <= lineBuffer_5141;
    end
    if (sel) begin
      lineBuffer_5143 <= lineBuffer_5142;
    end
    if (sel) begin
      lineBuffer_5144 <= lineBuffer_5143;
    end
    if (sel) begin
      lineBuffer_5145 <= lineBuffer_5144;
    end
    if (sel) begin
      lineBuffer_5146 <= lineBuffer_5145;
    end
    if (sel) begin
      lineBuffer_5147 <= lineBuffer_5146;
    end
    if (sel) begin
      lineBuffer_5148 <= lineBuffer_5147;
    end
    if (sel) begin
      lineBuffer_5149 <= lineBuffer_5148;
    end
    if (sel) begin
      lineBuffer_5150 <= lineBuffer_5149;
    end
    if (sel) begin
      lineBuffer_5151 <= lineBuffer_5150;
    end
    if (sel) begin
      lineBuffer_5152 <= lineBuffer_5151;
    end
    if (sel) begin
      lineBuffer_5153 <= lineBuffer_5152;
    end
    if (sel) begin
      lineBuffer_5154 <= lineBuffer_5153;
    end
    if (sel) begin
      lineBuffer_5155 <= lineBuffer_5154;
    end
    if (sel) begin
      lineBuffer_5156 <= lineBuffer_5155;
    end
    if (sel) begin
      lineBuffer_5157 <= lineBuffer_5156;
    end
    if (sel) begin
      lineBuffer_5158 <= lineBuffer_5157;
    end
    if (sel) begin
      lineBuffer_5159 <= lineBuffer_5158;
    end
    if (sel) begin
      lineBuffer_5160 <= lineBuffer_5159;
    end
    if (sel) begin
      lineBuffer_5161 <= lineBuffer_5160;
    end
    if (sel) begin
      lineBuffer_5162 <= lineBuffer_5161;
    end
    if (sel) begin
      lineBuffer_5163 <= lineBuffer_5162;
    end
    if (sel) begin
      lineBuffer_5164 <= lineBuffer_5163;
    end
    if (sel) begin
      lineBuffer_5165 <= lineBuffer_5164;
    end
    if (sel) begin
      lineBuffer_5166 <= lineBuffer_5165;
    end
    if (sel) begin
      lineBuffer_5167 <= lineBuffer_5166;
    end
    if (sel) begin
      lineBuffer_5168 <= lineBuffer_5167;
    end
    if (sel) begin
      lineBuffer_5169 <= lineBuffer_5168;
    end
    if (sel) begin
      lineBuffer_5170 <= lineBuffer_5169;
    end
    if (sel) begin
      lineBuffer_5171 <= lineBuffer_5170;
    end
    if (sel) begin
      lineBuffer_5172 <= lineBuffer_5171;
    end
    if (sel) begin
      lineBuffer_5173 <= lineBuffer_5172;
    end
    if (sel) begin
      lineBuffer_5174 <= lineBuffer_5173;
    end
    if (sel) begin
      lineBuffer_5175 <= lineBuffer_5174;
    end
    if (sel) begin
      lineBuffer_5176 <= lineBuffer_5175;
    end
    if (sel) begin
      lineBuffer_5177 <= lineBuffer_5176;
    end
    if (sel) begin
      lineBuffer_5178 <= lineBuffer_5177;
    end
    if (sel) begin
      lineBuffer_5179 <= lineBuffer_5178;
    end
    if (sel) begin
      lineBuffer_5180 <= lineBuffer_5179;
    end
    if (sel) begin
      lineBuffer_5181 <= lineBuffer_5180;
    end
    if (sel) begin
      lineBuffer_5182 <= lineBuffer_5181;
    end
    if (sel) begin
      lineBuffer_5183 <= lineBuffer_5182;
    end
    if (sel) begin
      lineBuffer_5184 <= lineBuffer_5183;
    end
    if (sel) begin
      lineBuffer_5185 <= lineBuffer_5184;
    end
    if (sel) begin
      lineBuffer_5186 <= lineBuffer_5185;
    end
    if (sel) begin
      lineBuffer_5187 <= lineBuffer_5186;
    end
    if (sel) begin
      lineBuffer_5188 <= lineBuffer_5187;
    end
    if (sel) begin
      lineBuffer_5189 <= lineBuffer_5188;
    end
    if (sel) begin
      lineBuffer_5190 <= lineBuffer_5189;
    end
    if (sel) begin
      lineBuffer_5191 <= lineBuffer_5190;
    end
    if (sel) begin
      lineBuffer_5192 <= lineBuffer_5191;
    end
    if (sel) begin
      lineBuffer_5193 <= lineBuffer_5192;
    end
    if (sel) begin
      lineBuffer_5194 <= lineBuffer_5193;
    end
    if (sel) begin
      lineBuffer_5195 <= lineBuffer_5194;
    end
    if (sel) begin
      lineBuffer_5196 <= lineBuffer_5195;
    end
    if (sel) begin
      lineBuffer_5197 <= lineBuffer_5196;
    end
    if (sel) begin
      lineBuffer_5198 <= lineBuffer_5197;
    end
    if (sel) begin
      lineBuffer_5199 <= lineBuffer_5198;
    end
    if (sel) begin
      lineBuffer_5200 <= lineBuffer_5199;
    end
    if (sel) begin
      lineBuffer_5201 <= lineBuffer_5200;
    end
    if (sel) begin
      lineBuffer_5202 <= lineBuffer_5201;
    end
    if (sel) begin
      lineBuffer_5203 <= lineBuffer_5202;
    end
    if (sel) begin
      lineBuffer_5204 <= lineBuffer_5203;
    end
    if (sel) begin
      lineBuffer_5205 <= lineBuffer_5204;
    end
    if (sel) begin
      lineBuffer_5206 <= lineBuffer_5205;
    end
    if (sel) begin
      lineBuffer_5207 <= lineBuffer_5206;
    end
    if (sel) begin
      lineBuffer_5208 <= lineBuffer_5207;
    end
    if (sel) begin
      lineBuffer_5209 <= lineBuffer_5208;
    end
    if (sel) begin
      lineBuffer_5210 <= lineBuffer_5209;
    end
    if (sel) begin
      lineBuffer_5211 <= lineBuffer_5210;
    end
    if (sel) begin
      lineBuffer_5212 <= lineBuffer_5211;
    end
    if (sel) begin
      lineBuffer_5213 <= lineBuffer_5212;
    end
    if (sel) begin
      lineBuffer_5214 <= lineBuffer_5213;
    end
    if (sel) begin
      lineBuffer_5215 <= lineBuffer_5214;
    end
    if (sel) begin
      lineBuffer_5216 <= lineBuffer_5215;
    end
    if (sel) begin
      lineBuffer_5217 <= lineBuffer_5216;
    end
    if (sel) begin
      lineBuffer_5218 <= lineBuffer_5217;
    end
    if (sel) begin
      lineBuffer_5219 <= lineBuffer_5218;
    end
    if (sel) begin
      lineBuffer_5220 <= lineBuffer_5219;
    end
    if (sel) begin
      lineBuffer_5221 <= lineBuffer_5220;
    end
    if (sel) begin
      lineBuffer_5222 <= lineBuffer_5221;
    end
    if (sel) begin
      lineBuffer_5223 <= lineBuffer_5222;
    end
    if (sel) begin
      lineBuffer_5224 <= lineBuffer_5223;
    end
    if (sel) begin
      lineBuffer_5225 <= lineBuffer_5224;
    end
    if (sel) begin
      lineBuffer_5226 <= lineBuffer_5225;
    end
    if (sel) begin
      lineBuffer_5227 <= lineBuffer_5226;
    end
    if (sel) begin
      lineBuffer_5228 <= lineBuffer_5227;
    end
    if (sel) begin
      lineBuffer_5229 <= lineBuffer_5228;
    end
    if (sel) begin
      lineBuffer_5230 <= lineBuffer_5229;
    end
    if (sel) begin
      lineBuffer_5231 <= lineBuffer_5230;
    end
    if (sel) begin
      lineBuffer_5232 <= lineBuffer_5231;
    end
    if (sel) begin
      lineBuffer_5233 <= lineBuffer_5232;
    end
    if (sel) begin
      lineBuffer_5234 <= lineBuffer_5233;
    end
    if (sel) begin
      lineBuffer_5235 <= lineBuffer_5234;
    end
    if (sel) begin
      lineBuffer_5236 <= lineBuffer_5235;
    end
    if (sel) begin
      lineBuffer_5237 <= lineBuffer_5236;
    end
    if (sel) begin
      lineBuffer_5238 <= lineBuffer_5237;
    end
    if (sel) begin
      lineBuffer_5239 <= lineBuffer_5238;
    end
    if (sel) begin
      lineBuffer_5240 <= lineBuffer_5239;
    end
    if (sel) begin
      lineBuffer_5241 <= lineBuffer_5240;
    end
    if (sel) begin
      lineBuffer_5242 <= lineBuffer_5241;
    end
    if (sel) begin
      lineBuffer_5243 <= lineBuffer_5242;
    end
    if (sel) begin
      lineBuffer_5244 <= lineBuffer_5243;
    end
    if (sel) begin
      lineBuffer_5245 <= lineBuffer_5244;
    end
    if (sel) begin
      lineBuffer_5246 <= lineBuffer_5245;
    end
    if (sel) begin
      lineBuffer_5247 <= lineBuffer_5246;
    end
    if (sel) begin
      lineBuffer_5248 <= lineBuffer_5247;
    end
    if (sel) begin
      lineBuffer_5249 <= lineBuffer_5248;
    end
    if (sel) begin
      lineBuffer_5250 <= lineBuffer_5249;
    end
    if (sel) begin
      lineBuffer_5251 <= lineBuffer_5250;
    end
    if (sel) begin
      lineBuffer_5252 <= lineBuffer_5251;
    end
    if (sel) begin
      lineBuffer_5253 <= lineBuffer_5252;
    end
    if (sel) begin
      lineBuffer_5254 <= lineBuffer_5253;
    end
    if (sel) begin
      lineBuffer_5255 <= lineBuffer_5254;
    end
    if (sel) begin
      lineBuffer_5256 <= lineBuffer_5255;
    end
    if (sel) begin
      lineBuffer_5257 <= lineBuffer_5256;
    end
    if (sel) begin
      lineBuffer_5258 <= lineBuffer_5257;
    end
    if (sel) begin
      lineBuffer_5259 <= lineBuffer_5258;
    end
    if (sel) begin
      lineBuffer_5260 <= lineBuffer_5259;
    end
    if (sel) begin
      lineBuffer_5261 <= lineBuffer_5260;
    end
    if (sel) begin
      lineBuffer_5262 <= lineBuffer_5261;
    end
    if (sel) begin
      lineBuffer_5263 <= lineBuffer_5262;
    end
    if (sel) begin
      lineBuffer_5264 <= lineBuffer_5263;
    end
    if (sel) begin
      lineBuffer_5265 <= lineBuffer_5264;
    end
    if (sel) begin
      lineBuffer_5266 <= lineBuffer_5265;
    end
    if (sel) begin
      lineBuffer_5267 <= lineBuffer_5266;
    end
    if (sel) begin
      lineBuffer_5268 <= lineBuffer_5267;
    end
    if (sel) begin
      lineBuffer_5269 <= lineBuffer_5268;
    end
    if (sel) begin
      lineBuffer_5270 <= lineBuffer_5269;
    end
    if (sel) begin
      lineBuffer_5271 <= lineBuffer_5270;
    end
    if (sel) begin
      lineBuffer_5272 <= lineBuffer_5271;
    end
    if (sel) begin
      lineBuffer_5273 <= lineBuffer_5272;
    end
    if (sel) begin
      lineBuffer_5274 <= lineBuffer_5273;
    end
    if (sel) begin
      lineBuffer_5275 <= lineBuffer_5274;
    end
    if (sel) begin
      lineBuffer_5276 <= lineBuffer_5275;
    end
    if (sel) begin
      lineBuffer_5277 <= lineBuffer_5276;
    end
    if (sel) begin
      lineBuffer_5278 <= lineBuffer_5277;
    end
    if (sel) begin
      lineBuffer_5279 <= lineBuffer_5278;
    end
    if (sel) begin
      lineBuffer_5280 <= lineBuffer_5279;
    end
    if (sel) begin
      lineBuffer_5281 <= lineBuffer_5280;
    end
    if (sel) begin
      lineBuffer_5282 <= lineBuffer_5281;
    end
    if (sel) begin
      lineBuffer_5283 <= lineBuffer_5282;
    end
    if (sel) begin
      lineBuffer_5284 <= lineBuffer_5283;
    end
    if (sel) begin
      lineBuffer_5285 <= lineBuffer_5284;
    end
    if (sel) begin
      lineBuffer_5286 <= lineBuffer_5285;
    end
    if (sel) begin
      lineBuffer_5287 <= lineBuffer_5286;
    end
    if (sel) begin
      lineBuffer_5288 <= lineBuffer_5287;
    end
    if (sel) begin
      lineBuffer_5289 <= lineBuffer_5288;
    end
    if (sel) begin
      lineBuffer_5290 <= lineBuffer_5289;
    end
    if (sel) begin
      lineBuffer_5291 <= lineBuffer_5290;
    end
    if (sel) begin
      lineBuffer_5292 <= lineBuffer_5291;
    end
    if (sel) begin
      lineBuffer_5293 <= lineBuffer_5292;
    end
    if (sel) begin
      lineBuffer_5294 <= lineBuffer_5293;
    end
    if (sel) begin
      lineBuffer_5295 <= lineBuffer_5294;
    end
    if (sel) begin
      lineBuffer_5296 <= lineBuffer_5295;
    end
    if (sel) begin
      lineBuffer_5297 <= lineBuffer_5296;
    end
    if (sel) begin
      lineBuffer_5298 <= lineBuffer_5297;
    end
    if (sel) begin
      lineBuffer_5299 <= lineBuffer_5298;
    end
    if (sel) begin
      lineBuffer_5300 <= lineBuffer_5299;
    end
    if (sel) begin
      lineBuffer_5301 <= lineBuffer_5300;
    end
    if (sel) begin
      lineBuffer_5302 <= lineBuffer_5301;
    end
    if (sel) begin
      lineBuffer_5303 <= lineBuffer_5302;
    end
    if (sel) begin
      lineBuffer_5304 <= lineBuffer_5303;
    end
    if (sel) begin
      lineBuffer_5305 <= lineBuffer_5304;
    end
    if (sel) begin
      lineBuffer_5306 <= lineBuffer_5305;
    end
    if (sel) begin
      lineBuffer_5307 <= lineBuffer_5306;
    end
    if (sel) begin
      lineBuffer_5308 <= lineBuffer_5307;
    end
    if (sel) begin
      lineBuffer_5309 <= lineBuffer_5308;
    end
    if (sel) begin
      lineBuffer_5310 <= lineBuffer_5309;
    end
    if (sel) begin
      lineBuffer_5311 <= lineBuffer_5310;
    end
    if (sel) begin
      lineBuffer_5312 <= lineBuffer_5311;
    end
    if (sel) begin
      lineBuffer_5313 <= lineBuffer_5312;
    end
    if (sel) begin
      lineBuffer_5314 <= lineBuffer_5313;
    end
    if (sel) begin
      lineBuffer_5315 <= lineBuffer_5314;
    end
    if (sel) begin
      lineBuffer_5316 <= lineBuffer_5315;
    end
    if (sel) begin
      lineBuffer_5317 <= lineBuffer_5316;
    end
    if (sel) begin
      lineBuffer_5318 <= lineBuffer_5317;
    end
    if (sel) begin
      lineBuffer_5319 <= lineBuffer_5318;
    end
    if (sel) begin
      lineBuffer_5320 <= lineBuffer_5319;
    end
    if (sel) begin
      lineBuffer_5321 <= lineBuffer_5320;
    end
    if (sel) begin
      lineBuffer_5322 <= lineBuffer_5321;
    end
    if (sel) begin
      lineBuffer_5323 <= lineBuffer_5322;
    end
    if (sel) begin
      lineBuffer_5324 <= lineBuffer_5323;
    end
    if (sel) begin
      lineBuffer_5325 <= lineBuffer_5324;
    end
    if (sel) begin
      lineBuffer_5326 <= lineBuffer_5325;
    end
    if (sel) begin
      lineBuffer_5327 <= lineBuffer_5326;
    end
    if (sel) begin
      lineBuffer_5328 <= lineBuffer_5327;
    end
    if (sel) begin
      lineBuffer_5329 <= lineBuffer_5328;
    end
    if (sel) begin
      lineBuffer_5330 <= lineBuffer_5329;
    end
    if (sel) begin
      lineBuffer_5331 <= lineBuffer_5330;
    end
    if (sel) begin
      lineBuffer_5332 <= lineBuffer_5331;
    end
    if (sel) begin
      lineBuffer_5333 <= lineBuffer_5332;
    end
    if (sel) begin
      lineBuffer_5334 <= lineBuffer_5333;
    end
    if (sel) begin
      lineBuffer_5335 <= lineBuffer_5334;
    end
    if (sel) begin
      lineBuffer_5336 <= lineBuffer_5335;
    end
    if (sel) begin
      lineBuffer_5337 <= lineBuffer_5336;
    end
    if (sel) begin
      lineBuffer_5338 <= lineBuffer_5337;
    end
    if (sel) begin
      lineBuffer_5339 <= lineBuffer_5338;
    end
    if (sel) begin
      lineBuffer_5340 <= lineBuffer_5339;
    end
    if (sel) begin
      lineBuffer_5341 <= lineBuffer_5340;
    end
    if (sel) begin
      lineBuffer_5342 <= lineBuffer_5341;
    end
    if (sel) begin
      lineBuffer_5343 <= lineBuffer_5342;
    end
    if (sel) begin
      lineBuffer_5344 <= lineBuffer_5343;
    end
    if (sel) begin
      lineBuffer_5345 <= lineBuffer_5344;
    end
    if (sel) begin
      lineBuffer_5346 <= lineBuffer_5345;
    end
    if (sel) begin
      lineBuffer_5347 <= lineBuffer_5346;
    end
    if (sel) begin
      lineBuffer_5348 <= lineBuffer_5347;
    end
    if (sel) begin
      lineBuffer_5349 <= lineBuffer_5348;
    end
    if (sel) begin
      lineBuffer_5350 <= lineBuffer_5349;
    end
    if (sel) begin
      lineBuffer_5351 <= lineBuffer_5350;
    end
    if (sel) begin
      lineBuffer_5352 <= lineBuffer_5351;
    end
    if (sel) begin
      lineBuffer_5353 <= lineBuffer_5352;
    end
    if (sel) begin
      lineBuffer_5354 <= lineBuffer_5353;
    end
    if (sel) begin
      lineBuffer_5355 <= lineBuffer_5354;
    end
    if (sel) begin
      lineBuffer_5356 <= lineBuffer_5355;
    end
    if (sel) begin
      lineBuffer_5357 <= lineBuffer_5356;
    end
    if (sel) begin
      lineBuffer_5358 <= lineBuffer_5357;
    end
    if (sel) begin
      lineBuffer_5359 <= lineBuffer_5358;
    end
    if (sel) begin
      lineBuffer_5360 <= lineBuffer_5359;
    end
    if (sel) begin
      lineBuffer_5361 <= lineBuffer_5360;
    end
    if (sel) begin
      lineBuffer_5362 <= lineBuffer_5361;
    end
    if (sel) begin
      lineBuffer_5363 <= lineBuffer_5362;
    end
    if (sel) begin
      lineBuffer_5364 <= lineBuffer_5363;
    end
    if (sel) begin
      lineBuffer_5365 <= lineBuffer_5364;
    end
    if (sel) begin
      lineBuffer_5366 <= lineBuffer_5365;
    end
    if (sel) begin
      lineBuffer_5367 <= lineBuffer_5366;
    end
    if (sel) begin
      lineBuffer_5368 <= lineBuffer_5367;
    end
    if (sel) begin
      lineBuffer_5369 <= lineBuffer_5368;
    end
    if (sel) begin
      lineBuffer_5370 <= lineBuffer_5369;
    end
    if (sel) begin
      lineBuffer_5371 <= lineBuffer_5370;
    end
    if (sel) begin
      lineBuffer_5372 <= lineBuffer_5371;
    end
    if (sel) begin
      lineBuffer_5373 <= lineBuffer_5372;
    end
    if (sel) begin
      lineBuffer_5374 <= lineBuffer_5373;
    end
    if (sel) begin
      lineBuffer_5375 <= lineBuffer_5374;
    end
    if (sel) begin
      lineBuffer_5376 <= lineBuffer_5375;
    end
    if (sel) begin
      lineBuffer_5377 <= lineBuffer_5376;
    end
    if (sel) begin
      lineBuffer_5378 <= lineBuffer_5377;
    end
    if (sel) begin
      lineBuffer_5379 <= lineBuffer_5378;
    end
    if (sel) begin
      lineBuffer_5380 <= lineBuffer_5379;
    end
    if (sel) begin
      lineBuffer_5381 <= lineBuffer_5380;
    end
    if (sel) begin
      lineBuffer_5382 <= lineBuffer_5381;
    end
    if (sel) begin
      lineBuffer_5383 <= lineBuffer_5382;
    end
    if (sel) begin
      lineBuffer_5384 <= lineBuffer_5383;
    end
    if (sel) begin
      lineBuffer_5385 <= lineBuffer_5384;
    end
    if (sel) begin
      lineBuffer_5386 <= lineBuffer_5385;
    end
    if (sel) begin
      lineBuffer_5387 <= lineBuffer_5386;
    end
    if (sel) begin
      lineBuffer_5388 <= lineBuffer_5387;
    end
    if (sel) begin
      lineBuffer_5389 <= lineBuffer_5388;
    end
    if (sel) begin
      lineBuffer_5390 <= lineBuffer_5389;
    end
    if (sel) begin
      lineBuffer_5391 <= lineBuffer_5390;
    end
    if (sel) begin
      lineBuffer_5392 <= lineBuffer_5391;
    end
    if (sel) begin
      lineBuffer_5393 <= lineBuffer_5392;
    end
    if (sel) begin
      lineBuffer_5394 <= lineBuffer_5393;
    end
    if (sel) begin
      lineBuffer_5395 <= lineBuffer_5394;
    end
    if (sel) begin
      lineBuffer_5396 <= lineBuffer_5395;
    end
    if (sel) begin
      lineBuffer_5397 <= lineBuffer_5396;
    end
    if (sel) begin
      lineBuffer_5398 <= lineBuffer_5397;
    end
    if (sel) begin
      lineBuffer_5399 <= lineBuffer_5398;
    end
    if (sel) begin
      lineBuffer_5400 <= lineBuffer_5399;
    end
    if (sel) begin
      lineBuffer_5401 <= lineBuffer_5400;
    end
    if (sel) begin
      lineBuffer_5402 <= lineBuffer_5401;
    end
    if (sel) begin
      lineBuffer_5403 <= lineBuffer_5402;
    end
    if (sel) begin
      lineBuffer_5404 <= lineBuffer_5403;
    end
    if (sel) begin
      lineBuffer_5405 <= lineBuffer_5404;
    end
    if (sel) begin
      lineBuffer_5406 <= lineBuffer_5405;
    end
    if (sel) begin
      lineBuffer_5407 <= lineBuffer_5406;
    end
    if (sel) begin
      lineBuffer_5408 <= lineBuffer_5407;
    end
    if (sel) begin
      lineBuffer_5409 <= lineBuffer_5408;
    end
    if (sel) begin
      lineBuffer_5410 <= lineBuffer_5409;
    end
    if (sel) begin
      lineBuffer_5411 <= lineBuffer_5410;
    end
    if (sel) begin
      lineBuffer_5412 <= lineBuffer_5411;
    end
    if (sel) begin
      lineBuffer_5413 <= lineBuffer_5412;
    end
    if (sel) begin
      lineBuffer_5414 <= lineBuffer_5413;
    end
    if (sel) begin
      lineBuffer_5415 <= lineBuffer_5414;
    end
    if (sel) begin
      lineBuffer_5416 <= lineBuffer_5415;
    end
    if (sel) begin
      lineBuffer_5417 <= lineBuffer_5416;
    end
    if (sel) begin
      lineBuffer_5418 <= lineBuffer_5417;
    end
    if (sel) begin
      lineBuffer_5419 <= lineBuffer_5418;
    end
    if (sel) begin
      lineBuffer_5420 <= lineBuffer_5419;
    end
    if (sel) begin
      lineBuffer_5421 <= lineBuffer_5420;
    end
    if (sel) begin
      lineBuffer_5422 <= lineBuffer_5421;
    end
    if (sel) begin
      lineBuffer_5423 <= lineBuffer_5422;
    end
    if (sel) begin
      lineBuffer_5424 <= lineBuffer_5423;
    end
    if (sel) begin
      lineBuffer_5425 <= lineBuffer_5424;
    end
    if (sel) begin
      lineBuffer_5426 <= lineBuffer_5425;
    end
    if (sel) begin
      lineBuffer_5427 <= lineBuffer_5426;
    end
    if (sel) begin
      lineBuffer_5428 <= lineBuffer_5427;
    end
    if (sel) begin
      lineBuffer_5429 <= lineBuffer_5428;
    end
    if (sel) begin
      lineBuffer_5430 <= lineBuffer_5429;
    end
    if (sel) begin
      lineBuffer_5431 <= lineBuffer_5430;
    end
    if (sel) begin
      lineBuffer_5432 <= lineBuffer_5431;
    end
    if (sel) begin
      lineBuffer_5433 <= lineBuffer_5432;
    end
    if (sel) begin
      lineBuffer_5434 <= lineBuffer_5433;
    end
    if (sel) begin
      lineBuffer_5435 <= lineBuffer_5434;
    end
    if (sel) begin
      lineBuffer_5436 <= lineBuffer_5435;
    end
    if (sel) begin
      lineBuffer_5437 <= lineBuffer_5436;
    end
    if (sel) begin
      lineBuffer_5438 <= lineBuffer_5437;
    end
    if (sel) begin
      lineBuffer_5439 <= lineBuffer_5438;
    end
    if (sel) begin
      lineBuffer_5440 <= lineBuffer_5439;
    end
    if (sel) begin
      lineBuffer_5441 <= lineBuffer_5440;
    end
    if (sel) begin
      lineBuffer_5442 <= lineBuffer_5441;
    end
    if (sel) begin
      lineBuffer_5443 <= lineBuffer_5442;
    end
    if (sel) begin
      lineBuffer_5444 <= lineBuffer_5443;
    end
    if (sel) begin
      lineBuffer_5445 <= lineBuffer_5444;
    end
    if (sel) begin
      lineBuffer_5446 <= lineBuffer_5445;
    end
    if (sel) begin
      lineBuffer_5447 <= lineBuffer_5446;
    end
    if (sel) begin
      lineBuffer_5448 <= lineBuffer_5447;
    end
    if (sel) begin
      lineBuffer_5449 <= lineBuffer_5448;
    end
    if (sel) begin
      lineBuffer_5450 <= lineBuffer_5449;
    end
    if (sel) begin
      lineBuffer_5451 <= lineBuffer_5450;
    end
    if (sel) begin
      lineBuffer_5452 <= lineBuffer_5451;
    end
    if (sel) begin
      lineBuffer_5453 <= lineBuffer_5452;
    end
    if (sel) begin
      lineBuffer_5454 <= lineBuffer_5453;
    end
    if (sel) begin
      lineBuffer_5455 <= lineBuffer_5454;
    end
    if (sel) begin
      lineBuffer_5456 <= lineBuffer_5455;
    end
    if (sel) begin
      lineBuffer_5457 <= lineBuffer_5456;
    end
    if (sel) begin
      lineBuffer_5458 <= lineBuffer_5457;
    end
    if (sel) begin
      lineBuffer_5459 <= lineBuffer_5458;
    end
    if (sel) begin
      lineBuffer_5460 <= lineBuffer_5459;
    end
    if (sel) begin
      lineBuffer_5461 <= lineBuffer_5460;
    end
    if (sel) begin
      lineBuffer_5462 <= lineBuffer_5461;
    end
    if (sel) begin
      lineBuffer_5463 <= lineBuffer_5462;
    end
    if (sel) begin
      lineBuffer_5464 <= lineBuffer_5463;
    end
    if (sel) begin
      lineBuffer_5465 <= lineBuffer_5464;
    end
    if (sel) begin
      lineBuffer_5466 <= lineBuffer_5465;
    end
    if (sel) begin
      lineBuffer_5467 <= lineBuffer_5466;
    end
    if (sel) begin
      lineBuffer_5468 <= lineBuffer_5467;
    end
    if (sel) begin
      lineBuffer_5469 <= lineBuffer_5468;
    end
    if (sel) begin
      lineBuffer_5470 <= lineBuffer_5469;
    end
    if (sel) begin
      lineBuffer_5471 <= lineBuffer_5470;
    end
    if (sel) begin
      lineBuffer_5472 <= lineBuffer_5471;
    end
    if (sel) begin
      lineBuffer_5473 <= lineBuffer_5472;
    end
    if (sel) begin
      lineBuffer_5474 <= lineBuffer_5473;
    end
    if (sel) begin
      lineBuffer_5475 <= lineBuffer_5474;
    end
    if (sel) begin
      lineBuffer_5476 <= lineBuffer_5475;
    end
    if (sel) begin
      lineBuffer_5477 <= lineBuffer_5476;
    end
    if (sel) begin
      lineBuffer_5478 <= lineBuffer_5477;
    end
    if (sel) begin
      lineBuffer_5479 <= lineBuffer_5478;
    end
    if (sel) begin
      lineBuffer_5480 <= lineBuffer_5479;
    end
    if (sel) begin
      lineBuffer_5481 <= lineBuffer_5480;
    end
    if (sel) begin
      lineBuffer_5482 <= lineBuffer_5481;
    end
    if (sel) begin
      lineBuffer_5483 <= lineBuffer_5482;
    end
    if (sel) begin
      lineBuffer_5484 <= lineBuffer_5483;
    end
    if (sel) begin
      lineBuffer_5485 <= lineBuffer_5484;
    end
    if (sel) begin
      lineBuffer_5486 <= lineBuffer_5485;
    end
    if (sel) begin
      lineBuffer_5487 <= lineBuffer_5486;
    end
    if (sel) begin
      lineBuffer_5488 <= lineBuffer_5487;
    end
    if (sel) begin
      lineBuffer_5489 <= lineBuffer_5488;
    end
    if (sel) begin
      lineBuffer_5490 <= lineBuffer_5489;
    end
    if (sel) begin
      lineBuffer_5491 <= lineBuffer_5490;
    end
    if (sel) begin
      lineBuffer_5492 <= lineBuffer_5491;
    end
    if (sel) begin
      lineBuffer_5493 <= lineBuffer_5492;
    end
    if (sel) begin
      lineBuffer_5494 <= lineBuffer_5493;
    end
    if (sel) begin
      lineBuffer_5495 <= lineBuffer_5494;
    end
    if (sel) begin
      lineBuffer_5496 <= lineBuffer_5495;
    end
    if (sel) begin
      lineBuffer_5497 <= lineBuffer_5496;
    end
    if (sel) begin
      lineBuffer_5498 <= lineBuffer_5497;
    end
    if (sel) begin
      lineBuffer_5499 <= lineBuffer_5498;
    end
    if (sel) begin
      lineBuffer_5500 <= lineBuffer_5499;
    end
    if (sel) begin
      lineBuffer_5501 <= lineBuffer_5500;
    end
    if (sel) begin
      lineBuffer_5502 <= lineBuffer_5501;
    end
    if (sel) begin
      lineBuffer_5503 <= lineBuffer_5502;
    end
    if (sel) begin
      lineBuffer_5504 <= lineBuffer_5503;
    end
    if (sel) begin
      lineBuffer_5505 <= lineBuffer_5504;
    end
    if (sel) begin
      lineBuffer_5506 <= lineBuffer_5505;
    end
    if (sel) begin
      lineBuffer_5507 <= lineBuffer_5506;
    end
    if (sel) begin
      lineBuffer_5508 <= lineBuffer_5507;
    end
    if (sel) begin
      lineBuffer_5509 <= lineBuffer_5508;
    end
    if (sel) begin
      lineBuffer_5510 <= lineBuffer_5509;
    end
    if (sel) begin
      lineBuffer_5511 <= lineBuffer_5510;
    end
    if (sel) begin
      lineBuffer_5512 <= lineBuffer_5511;
    end
    if (sel) begin
      lineBuffer_5513 <= lineBuffer_5512;
    end
    if (sel) begin
      lineBuffer_5514 <= lineBuffer_5513;
    end
    if (sel) begin
      lineBuffer_5515 <= lineBuffer_5514;
    end
    if (sel) begin
      lineBuffer_5516 <= lineBuffer_5515;
    end
    if (sel) begin
      lineBuffer_5517 <= lineBuffer_5516;
    end
    if (sel) begin
      lineBuffer_5518 <= lineBuffer_5517;
    end
    if (sel) begin
      lineBuffer_5519 <= lineBuffer_5518;
    end
    if (sel) begin
      lineBuffer_5520 <= lineBuffer_5519;
    end
    if (sel) begin
      lineBuffer_5521 <= lineBuffer_5520;
    end
    if (sel) begin
      lineBuffer_5522 <= lineBuffer_5521;
    end
    if (sel) begin
      lineBuffer_5523 <= lineBuffer_5522;
    end
    if (sel) begin
      lineBuffer_5524 <= lineBuffer_5523;
    end
    if (sel) begin
      lineBuffer_5525 <= lineBuffer_5524;
    end
    if (sel) begin
      lineBuffer_5526 <= lineBuffer_5525;
    end
    if (sel) begin
      lineBuffer_5527 <= lineBuffer_5526;
    end
    if (sel) begin
      lineBuffer_5528 <= lineBuffer_5527;
    end
    if (sel) begin
      lineBuffer_5529 <= lineBuffer_5528;
    end
    if (sel) begin
      lineBuffer_5530 <= lineBuffer_5529;
    end
    if (sel) begin
      lineBuffer_5531 <= lineBuffer_5530;
    end
    if (sel) begin
      lineBuffer_5532 <= lineBuffer_5531;
    end
    if (sel) begin
      lineBuffer_5533 <= lineBuffer_5532;
    end
    if (sel) begin
      lineBuffer_5534 <= lineBuffer_5533;
    end
    if (sel) begin
      lineBuffer_5535 <= lineBuffer_5534;
    end
    if (sel) begin
      lineBuffer_5536 <= lineBuffer_5535;
    end
    if (sel) begin
      lineBuffer_5537 <= lineBuffer_5536;
    end
    if (sel) begin
      lineBuffer_5538 <= lineBuffer_5537;
    end
    if (sel) begin
      lineBuffer_5539 <= lineBuffer_5538;
    end
    if (sel) begin
      lineBuffer_5540 <= lineBuffer_5539;
    end
    if (sel) begin
      lineBuffer_5541 <= lineBuffer_5540;
    end
    if (sel) begin
      lineBuffer_5542 <= lineBuffer_5541;
    end
    if (sel) begin
      lineBuffer_5543 <= lineBuffer_5542;
    end
    if (sel) begin
      lineBuffer_5544 <= lineBuffer_5543;
    end
    if (sel) begin
      lineBuffer_5545 <= lineBuffer_5544;
    end
    if (sel) begin
      lineBuffer_5546 <= lineBuffer_5545;
    end
    if (sel) begin
      lineBuffer_5547 <= lineBuffer_5546;
    end
    if (sel) begin
      lineBuffer_5548 <= lineBuffer_5547;
    end
    if (sel) begin
      lineBuffer_5549 <= lineBuffer_5548;
    end
    if (sel) begin
      lineBuffer_5550 <= lineBuffer_5549;
    end
    if (sel) begin
      lineBuffer_5551 <= lineBuffer_5550;
    end
    if (sel) begin
      lineBuffer_5552 <= lineBuffer_5551;
    end
    if (sel) begin
      lineBuffer_5553 <= lineBuffer_5552;
    end
    if (sel) begin
      lineBuffer_5554 <= lineBuffer_5553;
    end
    if (sel) begin
      lineBuffer_5555 <= lineBuffer_5554;
    end
    if (sel) begin
      lineBuffer_5556 <= lineBuffer_5555;
    end
    if (sel) begin
      lineBuffer_5557 <= lineBuffer_5556;
    end
    if (sel) begin
      lineBuffer_5558 <= lineBuffer_5557;
    end
    if (sel) begin
      lineBuffer_5559 <= lineBuffer_5558;
    end
    if (sel) begin
      lineBuffer_5560 <= lineBuffer_5559;
    end
    if (sel) begin
      lineBuffer_5561 <= lineBuffer_5560;
    end
    if (sel) begin
      lineBuffer_5562 <= lineBuffer_5561;
    end
    if (sel) begin
      lineBuffer_5563 <= lineBuffer_5562;
    end
    if (sel) begin
      lineBuffer_5564 <= lineBuffer_5563;
    end
    if (sel) begin
      lineBuffer_5565 <= lineBuffer_5564;
    end
    if (sel) begin
      lineBuffer_5566 <= lineBuffer_5565;
    end
    if (sel) begin
      lineBuffer_5567 <= lineBuffer_5566;
    end
    if (sel) begin
      lineBuffer_5568 <= lineBuffer_5567;
    end
    if (sel) begin
      lineBuffer_5569 <= lineBuffer_5568;
    end
    if (sel) begin
      lineBuffer_5570 <= lineBuffer_5569;
    end
    if (sel) begin
      lineBuffer_5571 <= lineBuffer_5570;
    end
    if (sel) begin
      lineBuffer_5572 <= lineBuffer_5571;
    end
    if (sel) begin
      lineBuffer_5573 <= lineBuffer_5572;
    end
    if (sel) begin
      lineBuffer_5574 <= lineBuffer_5573;
    end
    if (sel) begin
      lineBuffer_5575 <= lineBuffer_5574;
    end
    if (sel) begin
      lineBuffer_5576 <= lineBuffer_5575;
    end
    if (sel) begin
      lineBuffer_5577 <= lineBuffer_5576;
    end
    if (sel) begin
      lineBuffer_5578 <= lineBuffer_5577;
    end
    if (sel) begin
      lineBuffer_5579 <= lineBuffer_5578;
    end
    if (sel) begin
      lineBuffer_5580 <= lineBuffer_5579;
    end
    if (sel) begin
      lineBuffer_5581 <= lineBuffer_5580;
    end
    if (sel) begin
      lineBuffer_5582 <= lineBuffer_5581;
    end
    if (sel) begin
      lineBuffer_5583 <= lineBuffer_5582;
    end
    if (sel) begin
      lineBuffer_5584 <= lineBuffer_5583;
    end
    if (sel) begin
      lineBuffer_5585 <= lineBuffer_5584;
    end
    if (sel) begin
      lineBuffer_5586 <= lineBuffer_5585;
    end
    if (sel) begin
      lineBuffer_5587 <= lineBuffer_5586;
    end
    if (sel) begin
      lineBuffer_5588 <= lineBuffer_5587;
    end
    if (sel) begin
      lineBuffer_5589 <= lineBuffer_5588;
    end
    if (sel) begin
      lineBuffer_5590 <= lineBuffer_5589;
    end
    if (sel) begin
      lineBuffer_5591 <= lineBuffer_5590;
    end
    if (sel) begin
      lineBuffer_5592 <= lineBuffer_5591;
    end
    if (sel) begin
      lineBuffer_5593 <= lineBuffer_5592;
    end
    if (sel) begin
      lineBuffer_5594 <= lineBuffer_5593;
    end
    if (sel) begin
      lineBuffer_5595 <= lineBuffer_5594;
    end
    if (sel) begin
      lineBuffer_5596 <= lineBuffer_5595;
    end
    if (sel) begin
      lineBuffer_5597 <= lineBuffer_5596;
    end
    if (sel) begin
      lineBuffer_5598 <= lineBuffer_5597;
    end
    if (sel) begin
      lineBuffer_5599 <= lineBuffer_5598;
    end
    if (sel) begin
      lineBuffer_5600 <= lineBuffer_5599;
    end
    if (sel) begin
      lineBuffer_5601 <= lineBuffer_5600;
    end
    if (sel) begin
      lineBuffer_5602 <= lineBuffer_5601;
    end
    if (sel) begin
      lineBuffer_5603 <= lineBuffer_5602;
    end
    if (sel) begin
      lineBuffer_5604 <= lineBuffer_5603;
    end
    if (sel) begin
      lineBuffer_5605 <= lineBuffer_5604;
    end
    if (sel) begin
      lineBuffer_5606 <= lineBuffer_5605;
    end
    if (sel) begin
      lineBuffer_5607 <= lineBuffer_5606;
    end
    if (sel) begin
      lineBuffer_5608 <= lineBuffer_5607;
    end
    if (sel) begin
      lineBuffer_5609 <= lineBuffer_5608;
    end
    if (sel) begin
      lineBuffer_5610 <= lineBuffer_5609;
    end
    if (sel) begin
      lineBuffer_5611 <= lineBuffer_5610;
    end
    if (sel) begin
      lineBuffer_5612 <= lineBuffer_5611;
    end
    if (sel) begin
      lineBuffer_5613 <= lineBuffer_5612;
    end
    if (sel) begin
      lineBuffer_5614 <= lineBuffer_5613;
    end
    if (sel) begin
      lineBuffer_5615 <= lineBuffer_5614;
    end
    if (sel) begin
      lineBuffer_5616 <= lineBuffer_5615;
    end
    if (sel) begin
      lineBuffer_5617 <= lineBuffer_5616;
    end
    if (sel) begin
      lineBuffer_5618 <= lineBuffer_5617;
    end
    if (sel) begin
      lineBuffer_5619 <= lineBuffer_5618;
    end
    if (sel) begin
      lineBuffer_5620 <= lineBuffer_5619;
    end
    if (sel) begin
      lineBuffer_5621 <= lineBuffer_5620;
    end
    if (sel) begin
      lineBuffer_5622 <= lineBuffer_5621;
    end
    if (sel) begin
      lineBuffer_5623 <= lineBuffer_5622;
    end
    if (sel) begin
      lineBuffer_5624 <= lineBuffer_5623;
    end
    if (sel) begin
      lineBuffer_5625 <= lineBuffer_5624;
    end
    if (sel) begin
      lineBuffer_5626 <= lineBuffer_5625;
    end
    if (sel) begin
      lineBuffer_5627 <= lineBuffer_5626;
    end
    if (sel) begin
      lineBuffer_5628 <= lineBuffer_5627;
    end
    if (sel) begin
      lineBuffer_5629 <= lineBuffer_5628;
    end
    if (sel) begin
      lineBuffer_5630 <= lineBuffer_5629;
    end
    if (sel) begin
      lineBuffer_5631 <= lineBuffer_5630;
    end
    if (sel) begin
      lineBuffer_5632 <= lineBuffer_5631;
    end
    if (sel) begin
      lineBuffer_5633 <= lineBuffer_5632;
    end
    if (sel) begin
      lineBuffer_5634 <= lineBuffer_5633;
    end
    if (sel) begin
      lineBuffer_5635 <= lineBuffer_5634;
    end
    if (sel) begin
      lineBuffer_5636 <= lineBuffer_5635;
    end
    if (sel) begin
      lineBuffer_5637 <= lineBuffer_5636;
    end
    if (sel) begin
      lineBuffer_5638 <= lineBuffer_5637;
    end
    if (sel) begin
      lineBuffer_5639 <= lineBuffer_5638;
    end
    if (sel) begin
      lineBuffer_5640 <= lineBuffer_5639;
    end
    if (sel) begin
      lineBuffer_5641 <= lineBuffer_5640;
    end
    if (sel) begin
      lineBuffer_5642 <= lineBuffer_5641;
    end
    if (sel) begin
      lineBuffer_5643 <= lineBuffer_5642;
    end
    if (sel) begin
      lineBuffer_5644 <= lineBuffer_5643;
    end
    if (sel) begin
      lineBuffer_5645 <= lineBuffer_5644;
    end
    if (sel) begin
      lineBuffer_5646 <= lineBuffer_5645;
    end
    if (sel) begin
      lineBuffer_5647 <= lineBuffer_5646;
    end
    if (sel) begin
      lineBuffer_5648 <= lineBuffer_5647;
    end
    if (sel) begin
      lineBuffer_5649 <= lineBuffer_5648;
    end
    if (sel) begin
      lineBuffer_5650 <= lineBuffer_5649;
    end
    if (sel) begin
      lineBuffer_5651 <= lineBuffer_5650;
    end
    if (sel) begin
      lineBuffer_5652 <= lineBuffer_5651;
    end
    if (sel) begin
      lineBuffer_5653 <= lineBuffer_5652;
    end
    if (sel) begin
      lineBuffer_5654 <= lineBuffer_5653;
    end
    if (sel) begin
      lineBuffer_5655 <= lineBuffer_5654;
    end
    if (sel) begin
      lineBuffer_5656 <= lineBuffer_5655;
    end
    if (sel) begin
      lineBuffer_5657 <= lineBuffer_5656;
    end
    if (sel) begin
      lineBuffer_5658 <= lineBuffer_5657;
    end
    if (sel) begin
      lineBuffer_5659 <= lineBuffer_5658;
    end
    if (sel) begin
      lineBuffer_5660 <= lineBuffer_5659;
    end
    if (sel) begin
      lineBuffer_5661 <= lineBuffer_5660;
    end
    if (sel) begin
      lineBuffer_5662 <= lineBuffer_5661;
    end
    if (sel) begin
      lineBuffer_5663 <= lineBuffer_5662;
    end
    if (sel) begin
      lineBuffer_5664 <= lineBuffer_5663;
    end
    if (sel) begin
      lineBuffer_5665 <= lineBuffer_5664;
    end
    if (sel) begin
      lineBuffer_5666 <= lineBuffer_5665;
    end
    if (sel) begin
      lineBuffer_5667 <= lineBuffer_5666;
    end
    if (sel) begin
      lineBuffer_5668 <= lineBuffer_5667;
    end
    if (sel) begin
      lineBuffer_5669 <= lineBuffer_5668;
    end
    if (sel) begin
      lineBuffer_5670 <= lineBuffer_5669;
    end
    if (sel) begin
      lineBuffer_5671 <= lineBuffer_5670;
    end
    if (sel) begin
      lineBuffer_5672 <= lineBuffer_5671;
    end
    if (sel) begin
      lineBuffer_5673 <= lineBuffer_5672;
    end
    if (sel) begin
      lineBuffer_5674 <= lineBuffer_5673;
    end
    if (sel) begin
      lineBuffer_5675 <= lineBuffer_5674;
    end
    if (sel) begin
      lineBuffer_5676 <= lineBuffer_5675;
    end
    if (sel) begin
      lineBuffer_5677 <= lineBuffer_5676;
    end
    if (sel) begin
      lineBuffer_5678 <= lineBuffer_5677;
    end
    if (sel) begin
      lineBuffer_5679 <= lineBuffer_5678;
    end
    if (sel) begin
      lineBuffer_5680 <= lineBuffer_5679;
    end
    if (sel) begin
      lineBuffer_5681 <= lineBuffer_5680;
    end
    if (sel) begin
      lineBuffer_5682 <= lineBuffer_5681;
    end
    if (sel) begin
      lineBuffer_5683 <= lineBuffer_5682;
    end
    if (sel) begin
      lineBuffer_5684 <= lineBuffer_5683;
    end
    if (sel) begin
      lineBuffer_5685 <= lineBuffer_5684;
    end
    if (sel) begin
      lineBuffer_5686 <= lineBuffer_5685;
    end
    if (sel) begin
      lineBuffer_5687 <= lineBuffer_5686;
    end
    if (sel) begin
      lineBuffer_5688 <= lineBuffer_5687;
    end
    if (sel) begin
      lineBuffer_5689 <= lineBuffer_5688;
    end
    if (sel) begin
      lineBuffer_5690 <= lineBuffer_5689;
    end
    if (sel) begin
      lineBuffer_5691 <= lineBuffer_5690;
    end
    if (sel) begin
      lineBuffer_5692 <= lineBuffer_5691;
    end
    if (sel) begin
      lineBuffer_5693 <= lineBuffer_5692;
    end
    if (sel) begin
      lineBuffer_5694 <= lineBuffer_5693;
    end
    if (sel) begin
      lineBuffer_5695 <= lineBuffer_5694;
    end
    if (sel) begin
      lineBuffer_5696 <= lineBuffer_5695;
    end
    if (sel) begin
      lineBuffer_5697 <= lineBuffer_5696;
    end
    if (sel) begin
      lineBuffer_5698 <= lineBuffer_5697;
    end
    if (sel) begin
      lineBuffer_5699 <= lineBuffer_5698;
    end
    if (sel) begin
      lineBuffer_5700 <= lineBuffer_5699;
    end
    if (sel) begin
      lineBuffer_5701 <= lineBuffer_5700;
    end
    if (sel) begin
      lineBuffer_5702 <= lineBuffer_5701;
    end
    if (sel) begin
      lineBuffer_5703 <= lineBuffer_5702;
    end
    if (sel) begin
      lineBuffer_5704 <= lineBuffer_5703;
    end
    if (sel) begin
      lineBuffer_5705 <= lineBuffer_5704;
    end
    if (sel) begin
      lineBuffer_5706 <= lineBuffer_5705;
    end
    if (sel) begin
      lineBuffer_5707 <= lineBuffer_5706;
    end
    if (sel) begin
      lineBuffer_5708 <= lineBuffer_5707;
    end
    if (sel) begin
      lineBuffer_5709 <= lineBuffer_5708;
    end
    if (sel) begin
      lineBuffer_5710 <= lineBuffer_5709;
    end
    if (sel) begin
      lineBuffer_5711 <= lineBuffer_5710;
    end
    if (sel) begin
      lineBuffer_5712 <= lineBuffer_5711;
    end
    if (sel) begin
      lineBuffer_5713 <= lineBuffer_5712;
    end
    if (sel) begin
      lineBuffer_5714 <= lineBuffer_5713;
    end
    if (sel) begin
      lineBuffer_5715 <= lineBuffer_5714;
    end
    if (sel) begin
      lineBuffer_5716 <= lineBuffer_5715;
    end
    if (sel) begin
      lineBuffer_5717 <= lineBuffer_5716;
    end
    if (sel) begin
      lineBuffer_5718 <= lineBuffer_5717;
    end
    if (sel) begin
      lineBuffer_5719 <= lineBuffer_5718;
    end
    if (sel) begin
      lineBuffer_5720 <= lineBuffer_5719;
    end
    if (sel) begin
      lineBuffer_5721 <= lineBuffer_5720;
    end
    if (sel) begin
      lineBuffer_5722 <= lineBuffer_5721;
    end
    if (sel) begin
      lineBuffer_5723 <= lineBuffer_5722;
    end
    if (sel) begin
      lineBuffer_5724 <= lineBuffer_5723;
    end
    if (sel) begin
      lineBuffer_5725 <= lineBuffer_5724;
    end
    if (sel) begin
      lineBuffer_5726 <= lineBuffer_5725;
    end
    if (sel) begin
      lineBuffer_5727 <= lineBuffer_5726;
    end
    if (sel) begin
      lineBuffer_5728 <= lineBuffer_5727;
    end
    if (sel) begin
      lineBuffer_5729 <= lineBuffer_5728;
    end
    if (sel) begin
      lineBuffer_5730 <= lineBuffer_5729;
    end
    if (sel) begin
      lineBuffer_5731 <= lineBuffer_5730;
    end
    if (sel) begin
      lineBuffer_5732 <= lineBuffer_5731;
    end
    if (sel) begin
      lineBuffer_5733 <= lineBuffer_5732;
    end
    if (sel) begin
      lineBuffer_5734 <= lineBuffer_5733;
    end
    if (sel) begin
      lineBuffer_5735 <= lineBuffer_5734;
    end
    if (sel) begin
      lineBuffer_5736 <= lineBuffer_5735;
    end
    if (sel) begin
      lineBuffer_5737 <= lineBuffer_5736;
    end
    if (sel) begin
      lineBuffer_5738 <= lineBuffer_5737;
    end
    if (sel) begin
      lineBuffer_5739 <= lineBuffer_5738;
    end
    if (sel) begin
      lineBuffer_5740 <= lineBuffer_5739;
    end
    if (sel) begin
      lineBuffer_5741 <= lineBuffer_5740;
    end
    if (sel) begin
      lineBuffer_5742 <= lineBuffer_5741;
    end
    if (sel) begin
      lineBuffer_5743 <= lineBuffer_5742;
    end
    if (sel) begin
      lineBuffer_5744 <= lineBuffer_5743;
    end
    if (sel) begin
      lineBuffer_5745 <= lineBuffer_5744;
    end
    if (sel) begin
      lineBuffer_5746 <= lineBuffer_5745;
    end
    if (sel) begin
      lineBuffer_5747 <= lineBuffer_5746;
    end
    if (sel) begin
      lineBuffer_5748 <= lineBuffer_5747;
    end
    if (sel) begin
      lineBuffer_5749 <= lineBuffer_5748;
    end
    if (sel) begin
      lineBuffer_5750 <= lineBuffer_5749;
    end
    if (sel) begin
      lineBuffer_5751 <= lineBuffer_5750;
    end
    if (sel) begin
      lineBuffer_5752 <= lineBuffer_5751;
    end
    if (sel) begin
      lineBuffer_5753 <= lineBuffer_5752;
    end
    if (sel) begin
      lineBuffer_5754 <= lineBuffer_5753;
    end
    if (sel) begin
      lineBuffer_5755 <= lineBuffer_5754;
    end
    if (sel) begin
      lineBuffer_5756 <= lineBuffer_5755;
    end
    if (sel) begin
      lineBuffer_5757 <= lineBuffer_5756;
    end
    if (sel) begin
      lineBuffer_5758 <= lineBuffer_5757;
    end
    if (sel) begin
      lineBuffer_5759 <= lineBuffer_5758;
    end
    if (sel) begin
      lineBuffer_5760 <= lineBuffer_5759;
    end
    if (sel) begin
      lineBuffer_5761 <= lineBuffer_5760;
    end
    if (sel) begin
      lineBuffer_5762 <= lineBuffer_5761;
    end
    if (sel) begin
      lineBuffer_5763 <= lineBuffer_5762;
    end
    if (sel) begin
      lineBuffer_5764 <= lineBuffer_5763;
    end
    if (sel) begin
      lineBuffer_5765 <= lineBuffer_5764;
    end
    if (sel) begin
      lineBuffer_5766 <= lineBuffer_5765;
    end
    if (sel) begin
      lineBuffer_5767 <= lineBuffer_5766;
    end
    if (sel) begin
      lineBuffer_5768 <= lineBuffer_5767;
    end
    if (sel) begin
      lineBuffer_5769 <= lineBuffer_5768;
    end
    if (sel) begin
      lineBuffer_5770 <= lineBuffer_5769;
    end
    if (sel) begin
      lineBuffer_5771 <= lineBuffer_5770;
    end
    if (sel) begin
      lineBuffer_5772 <= lineBuffer_5771;
    end
    if (sel) begin
      lineBuffer_5773 <= lineBuffer_5772;
    end
    if (sel) begin
      lineBuffer_5774 <= lineBuffer_5773;
    end
    if (sel) begin
      lineBuffer_5775 <= lineBuffer_5774;
    end
    if (sel) begin
      lineBuffer_5776 <= lineBuffer_5775;
    end
    if (sel) begin
      lineBuffer_5777 <= lineBuffer_5776;
    end
    if (sel) begin
      lineBuffer_5778 <= lineBuffer_5777;
    end
    if (sel) begin
      lineBuffer_5779 <= lineBuffer_5778;
    end
    if (sel) begin
      lineBuffer_5780 <= lineBuffer_5779;
    end
    if (sel) begin
      lineBuffer_5781 <= lineBuffer_5780;
    end
    if (sel) begin
      lineBuffer_5782 <= lineBuffer_5781;
    end
    if (sel) begin
      lineBuffer_5783 <= lineBuffer_5782;
    end
    if (sel) begin
      lineBuffer_5784 <= lineBuffer_5783;
    end
    if (sel) begin
      lineBuffer_5785 <= lineBuffer_5784;
    end
    if (sel) begin
      lineBuffer_5786 <= lineBuffer_5785;
    end
    if (sel) begin
      lineBuffer_5787 <= lineBuffer_5786;
    end
    if (sel) begin
      lineBuffer_5788 <= lineBuffer_5787;
    end
    if (sel) begin
      lineBuffer_5789 <= lineBuffer_5788;
    end
    if (sel) begin
      lineBuffer_5790 <= lineBuffer_5789;
    end
    if (sel) begin
      lineBuffer_5791 <= lineBuffer_5790;
    end
    if (sel) begin
      lineBuffer_5792 <= lineBuffer_5791;
    end
    if (sel) begin
      lineBuffer_5793 <= lineBuffer_5792;
    end
    if (sel) begin
      lineBuffer_5794 <= lineBuffer_5793;
    end
    if (sel) begin
      lineBuffer_5795 <= lineBuffer_5794;
    end
    if (sel) begin
      lineBuffer_5796 <= lineBuffer_5795;
    end
    if (sel) begin
      lineBuffer_5797 <= lineBuffer_5796;
    end
    if (sel) begin
      lineBuffer_5798 <= lineBuffer_5797;
    end
    if (sel) begin
      lineBuffer_5799 <= lineBuffer_5798;
    end
    if (sel) begin
      lineBuffer_5800 <= lineBuffer_5799;
    end
    if (sel) begin
      lineBuffer_5801 <= lineBuffer_5800;
    end
    if (sel) begin
      lineBuffer_5802 <= lineBuffer_5801;
    end
    if (sel) begin
      lineBuffer_5803 <= lineBuffer_5802;
    end
    if (sel) begin
      lineBuffer_5804 <= lineBuffer_5803;
    end
    if (sel) begin
      lineBuffer_5805 <= lineBuffer_5804;
    end
    if (sel) begin
      lineBuffer_5806 <= lineBuffer_5805;
    end
    if (sel) begin
      lineBuffer_5807 <= lineBuffer_5806;
    end
    if (sel) begin
      lineBuffer_5808 <= lineBuffer_5807;
    end
    if (sel) begin
      lineBuffer_5809 <= lineBuffer_5808;
    end
    if (sel) begin
      lineBuffer_5810 <= lineBuffer_5809;
    end
    if (sel) begin
      lineBuffer_5811 <= lineBuffer_5810;
    end
    if (sel) begin
      lineBuffer_5812 <= lineBuffer_5811;
    end
    if (sel) begin
      lineBuffer_5813 <= lineBuffer_5812;
    end
    if (sel) begin
      lineBuffer_5814 <= lineBuffer_5813;
    end
    if (sel) begin
      lineBuffer_5815 <= lineBuffer_5814;
    end
    if (sel) begin
      lineBuffer_5816 <= lineBuffer_5815;
    end
    if (sel) begin
      lineBuffer_5817 <= lineBuffer_5816;
    end
    if (sel) begin
      lineBuffer_5818 <= lineBuffer_5817;
    end
    if (sel) begin
      lineBuffer_5819 <= lineBuffer_5818;
    end
    if (sel) begin
      lineBuffer_5820 <= lineBuffer_5819;
    end
    if (sel) begin
      lineBuffer_5821 <= lineBuffer_5820;
    end
    if (sel) begin
      lineBuffer_5822 <= lineBuffer_5821;
    end
    if (sel) begin
      lineBuffer_5823 <= lineBuffer_5822;
    end
    if (sel) begin
      lineBuffer_5824 <= lineBuffer_5823;
    end
    if (sel) begin
      lineBuffer_5825 <= lineBuffer_5824;
    end
    if (sel) begin
      lineBuffer_5826 <= lineBuffer_5825;
    end
    if (sel) begin
      lineBuffer_5827 <= lineBuffer_5826;
    end
    if (sel) begin
      lineBuffer_5828 <= lineBuffer_5827;
    end
    if (sel) begin
      lineBuffer_5829 <= lineBuffer_5828;
    end
    if (sel) begin
      lineBuffer_5830 <= lineBuffer_5829;
    end
    if (sel) begin
      lineBuffer_5831 <= lineBuffer_5830;
    end
    if (sel) begin
      lineBuffer_5832 <= lineBuffer_5831;
    end
    if (sel) begin
      lineBuffer_5833 <= lineBuffer_5832;
    end
    if (sel) begin
      lineBuffer_5834 <= lineBuffer_5833;
    end
    if (sel) begin
      lineBuffer_5835 <= lineBuffer_5834;
    end
    if (sel) begin
      lineBuffer_5836 <= lineBuffer_5835;
    end
    if (sel) begin
      lineBuffer_5837 <= lineBuffer_5836;
    end
    if (sel) begin
      lineBuffer_5838 <= lineBuffer_5837;
    end
    if (sel) begin
      lineBuffer_5839 <= lineBuffer_5838;
    end
    if (sel) begin
      lineBuffer_5840 <= lineBuffer_5839;
    end
    if (sel) begin
      lineBuffer_5841 <= lineBuffer_5840;
    end
    if (sel) begin
      lineBuffer_5842 <= lineBuffer_5841;
    end
    if (sel) begin
      lineBuffer_5843 <= lineBuffer_5842;
    end
    if (sel) begin
      lineBuffer_5844 <= lineBuffer_5843;
    end
    if (sel) begin
      lineBuffer_5845 <= lineBuffer_5844;
    end
    if (sel) begin
      lineBuffer_5846 <= lineBuffer_5845;
    end
    if (sel) begin
      lineBuffer_5847 <= lineBuffer_5846;
    end
    if (sel) begin
      lineBuffer_5848 <= lineBuffer_5847;
    end
    if (sel) begin
      lineBuffer_5849 <= lineBuffer_5848;
    end
    if (sel) begin
      lineBuffer_5850 <= lineBuffer_5849;
    end
    if (sel) begin
      lineBuffer_5851 <= lineBuffer_5850;
    end
    if (sel) begin
      lineBuffer_5852 <= lineBuffer_5851;
    end
    if (sel) begin
      lineBuffer_5853 <= lineBuffer_5852;
    end
    if (sel) begin
      lineBuffer_5854 <= lineBuffer_5853;
    end
    if (sel) begin
      lineBuffer_5855 <= lineBuffer_5854;
    end
    if (sel) begin
      lineBuffer_5856 <= lineBuffer_5855;
    end
    if (sel) begin
      lineBuffer_5857 <= lineBuffer_5856;
    end
    if (sel) begin
      lineBuffer_5858 <= lineBuffer_5857;
    end
    if (sel) begin
      lineBuffer_5859 <= lineBuffer_5858;
    end
    if (sel) begin
      lineBuffer_5860 <= lineBuffer_5859;
    end
    if (sel) begin
      lineBuffer_5861 <= lineBuffer_5860;
    end
    if (sel) begin
      lineBuffer_5862 <= lineBuffer_5861;
    end
    if (sel) begin
      lineBuffer_5863 <= lineBuffer_5862;
    end
    if (sel) begin
      lineBuffer_5864 <= lineBuffer_5863;
    end
    if (sel) begin
      lineBuffer_5865 <= lineBuffer_5864;
    end
    if (sel) begin
      lineBuffer_5866 <= lineBuffer_5865;
    end
    if (sel) begin
      lineBuffer_5867 <= lineBuffer_5866;
    end
    if (sel) begin
      lineBuffer_5868 <= lineBuffer_5867;
    end
    if (sel) begin
      lineBuffer_5869 <= lineBuffer_5868;
    end
    if (sel) begin
      lineBuffer_5870 <= lineBuffer_5869;
    end
    if (sel) begin
      lineBuffer_5871 <= lineBuffer_5870;
    end
    if (sel) begin
      lineBuffer_5872 <= lineBuffer_5871;
    end
    if (sel) begin
      lineBuffer_5873 <= lineBuffer_5872;
    end
    if (sel) begin
      lineBuffer_5874 <= lineBuffer_5873;
    end
    if (sel) begin
      lineBuffer_5875 <= lineBuffer_5874;
    end
    if (sel) begin
      lineBuffer_5876 <= lineBuffer_5875;
    end
    if (sel) begin
      lineBuffer_5877 <= lineBuffer_5876;
    end
    if (sel) begin
      lineBuffer_5878 <= lineBuffer_5877;
    end
    if (sel) begin
      lineBuffer_5879 <= lineBuffer_5878;
    end
    if (sel) begin
      lineBuffer_5880 <= lineBuffer_5879;
    end
    if (sel) begin
      lineBuffer_5881 <= lineBuffer_5880;
    end
    if (sel) begin
      lineBuffer_5882 <= lineBuffer_5881;
    end
    if (sel) begin
      lineBuffer_5883 <= lineBuffer_5882;
    end
    if (sel) begin
      lineBuffer_5884 <= lineBuffer_5883;
    end
    if (sel) begin
      lineBuffer_5885 <= lineBuffer_5884;
    end
    if (sel) begin
      lineBuffer_5886 <= lineBuffer_5885;
    end
    if (sel) begin
      lineBuffer_5887 <= lineBuffer_5886;
    end
    if (sel) begin
      lineBuffer_5888 <= lineBuffer_5887;
    end
    if (sel) begin
      lineBuffer_5889 <= lineBuffer_5888;
    end
    if (sel) begin
      lineBuffer_5890 <= lineBuffer_5889;
    end
    if (sel) begin
      lineBuffer_5891 <= lineBuffer_5890;
    end
    if (sel) begin
      lineBuffer_5892 <= lineBuffer_5891;
    end
    if (sel) begin
      lineBuffer_5893 <= lineBuffer_5892;
    end
    if (sel) begin
      lineBuffer_5894 <= lineBuffer_5893;
    end
    if (sel) begin
      lineBuffer_5895 <= lineBuffer_5894;
    end
    if (sel) begin
      lineBuffer_5896 <= lineBuffer_5895;
    end
    if (sel) begin
      lineBuffer_5897 <= lineBuffer_5896;
    end
    if (sel) begin
      lineBuffer_5898 <= lineBuffer_5897;
    end
    if (sel) begin
      lineBuffer_5899 <= lineBuffer_5898;
    end
    if (sel) begin
      lineBuffer_5900 <= lineBuffer_5899;
    end
    if (sel) begin
      lineBuffer_5901 <= lineBuffer_5900;
    end
    if (sel) begin
      lineBuffer_5902 <= lineBuffer_5901;
    end
    if (sel) begin
      lineBuffer_5903 <= lineBuffer_5902;
    end
    if (sel) begin
      lineBuffer_5904 <= lineBuffer_5903;
    end
    if (sel) begin
      lineBuffer_5905 <= lineBuffer_5904;
    end
    if (sel) begin
      lineBuffer_5906 <= lineBuffer_5905;
    end
    if (sel) begin
      lineBuffer_5907 <= lineBuffer_5906;
    end
    if (sel) begin
      lineBuffer_5908 <= lineBuffer_5907;
    end
    if (sel) begin
      lineBuffer_5909 <= lineBuffer_5908;
    end
    if (sel) begin
      lineBuffer_5910 <= lineBuffer_5909;
    end
    if (sel) begin
      lineBuffer_5911 <= lineBuffer_5910;
    end
    if (sel) begin
      lineBuffer_5912 <= lineBuffer_5911;
    end
    if (sel) begin
      lineBuffer_5913 <= lineBuffer_5912;
    end
    if (sel) begin
      lineBuffer_5914 <= lineBuffer_5913;
    end
    if (sel) begin
      lineBuffer_5915 <= lineBuffer_5914;
    end
    if (sel) begin
      lineBuffer_5916 <= lineBuffer_5915;
    end
    if (sel) begin
      lineBuffer_5917 <= lineBuffer_5916;
    end
    if (sel) begin
      lineBuffer_5918 <= lineBuffer_5917;
    end
    if (sel) begin
      lineBuffer_5919 <= lineBuffer_5918;
    end
    if (sel) begin
      lineBuffer_5920 <= lineBuffer_5919;
    end
    if (sel) begin
      lineBuffer_5921 <= lineBuffer_5920;
    end
    if (sel) begin
      lineBuffer_5922 <= lineBuffer_5921;
    end
    if (sel) begin
      lineBuffer_5923 <= lineBuffer_5922;
    end
    if (sel) begin
      lineBuffer_5924 <= lineBuffer_5923;
    end
    if (sel) begin
      lineBuffer_5925 <= lineBuffer_5924;
    end
    if (sel) begin
      lineBuffer_5926 <= lineBuffer_5925;
    end
    if (sel) begin
      lineBuffer_5927 <= lineBuffer_5926;
    end
    if (sel) begin
      lineBuffer_5928 <= lineBuffer_5927;
    end
    if (sel) begin
      lineBuffer_5929 <= lineBuffer_5928;
    end
    if (sel) begin
      lineBuffer_5930 <= lineBuffer_5929;
    end
    if (sel) begin
      lineBuffer_5931 <= lineBuffer_5930;
    end
    if (sel) begin
      lineBuffer_5932 <= lineBuffer_5931;
    end
    if (sel) begin
      lineBuffer_5933 <= lineBuffer_5932;
    end
    if (sel) begin
      lineBuffer_5934 <= lineBuffer_5933;
    end
    if (sel) begin
      lineBuffer_5935 <= lineBuffer_5934;
    end
    if (sel) begin
      lineBuffer_5936 <= lineBuffer_5935;
    end
    if (sel) begin
      lineBuffer_5937 <= lineBuffer_5936;
    end
    if (sel) begin
      lineBuffer_5938 <= lineBuffer_5937;
    end
    if (sel) begin
      lineBuffer_5939 <= lineBuffer_5938;
    end
    if (sel) begin
      lineBuffer_5940 <= lineBuffer_5939;
    end
    if (sel) begin
      lineBuffer_5941 <= lineBuffer_5940;
    end
    if (sel) begin
      lineBuffer_5942 <= lineBuffer_5941;
    end
    if (sel) begin
      lineBuffer_5943 <= lineBuffer_5942;
    end
    if (sel) begin
      lineBuffer_5944 <= lineBuffer_5943;
    end
    if (sel) begin
      lineBuffer_5945 <= lineBuffer_5944;
    end
    if (sel) begin
      lineBuffer_5946 <= lineBuffer_5945;
    end
    if (sel) begin
      lineBuffer_5947 <= lineBuffer_5946;
    end
    if (sel) begin
      lineBuffer_5948 <= lineBuffer_5947;
    end
    if (sel) begin
      lineBuffer_5949 <= lineBuffer_5948;
    end
    if (sel) begin
      lineBuffer_5950 <= lineBuffer_5949;
    end
    if (sel) begin
      lineBuffer_5951 <= lineBuffer_5950;
    end
    if (sel) begin
      lineBuffer_5952 <= lineBuffer_5951;
    end
    if (sel) begin
      lineBuffer_5953 <= lineBuffer_5952;
    end
    if (sel) begin
      lineBuffer_5954 <= lineBuffer_5953;
    end
    if (sel) begin
      lineBuffer_5955 <= lineBuffer_5954;
    end
    if (sel) begin
      lineBuffer_5956 <= lineBuffer_5955;
    end
    if (sel) begin
      lineBuffer_5957 <= lineBuffer_5956;
    end
    if (sel) begin
      lineBuffer_5958 <= lineBuffer_5957;
    end
    if (sel) begin
      lineBuffer_5959 <= lineBuffer_5958;
    end
    if (sel) begin
      lineBuffer_5960 <= lineBuffer_5959;
    end
    if (sel) begin
      lineBuffer_5961 <= lineBuffer_5960;
    end
    if (sel) begin
      lineBuffer_5962 <= lineBuffer_5961;
    end
    if (sel) begin
      lineBuffer_5963 <= lineBuffer_5962;
    end
    if (sel) begin
      lineBuffer_5964 <= lineBuffer_5963;
    end
    if (sel) begin
      lineBuffer_5965 <= lineBuffer_5964;
    end
    if (sel) begin
      lineBuffer_5966 <= lineBuffer_5965;
    end
    if (sel) begin
      lineBuffer_5967 <= lineBuffer_5966;
    end
    if (sel) begin
      lineBuffer_5968 <= lineBuffer_5967;
    end
    if (sel) begin
      lineBuffer_5969 <= lineBuffer_5968;
    end
    if (sel) begin
      lineBuffer_5970 <= lineBuffer_5969;
    end
    if (sel) begin
      lineBuffer_5971 <= lineBuffer_5970;
    end
    if (sel) begin
      lineBuffer_5972 <= lineBuffer_5971;
    end
    if (sel) begin
      lineBuffer_5973 <= lineBuffer_5972;
    end
    if (sel) begin
      lineBuffer_5974 <= lineBuffer_5973;
    end
    if (sel) begin
      lineBuffer_5975 <= lineBuffer_5974;
    end
    if (sel) begin
      lineBuffer_5976 <= lineBuffer_5975;
    end
    if (sel) begin
      lineBuffer_5977 <= lineBuffer_5976;
    end
    if (sel) begin
      lineBuffer_5978 <= lineBuffer_5977;
    end
    if (sel) begin
      lineBuffer_5979 <= lineBuffer_5978;
    end
    if (sel) begin
      lineBuffer_5980 <= lineBuffer_5979;
    end
    if (sel) begin
      lineBuffer_5981 <= lineBuffer_5980;
    end
    if (sel) begin
      lineBuffer_5982 <= lineBuffer_5981;
    end
    if (sel) begin
      lineBuffer_5983 <= lineBuffer_5982;
    end
    if (sel) begin
      lineBuffer_5984 <= lineBuffer_5983;
    end
    if (sel) begin
      lineBuffer_5985 <= lineBuffer_5984;
    end
    if (sel) begin
      lineBuffer_5986 <= lineBuffer_5985;
    end
    if (sel) begin
      lineBuffer_5987 <= lineBuffer_5986;
    end
    if (sel) begin
      lineBuffer_5988 <= lineBuffer_5987;
    end
    if (sel) begin
      lineBuffer_5989 <= lineBuffer_5988;
    end
    if (sel) begin
      lineBuffer_5990 <= lineBuffer_5989;
    end
    if (sel) begin
      lineBuffer_5991 <= lineBuffer_5990;
    end
    if (sel) begin
      lineBuffer_5992 <= lineBuffer_5991;
    end
    if (sel) begin
      lineBuffer_5993 <= lineBuffer_5992;
    end
    if (sel) begin
      lineBuffer_5994 <= lineBuffer_5993;
    end
    if (sel) begin
      lineBuffer_5995 <= lineBuffer_5994;
    end
    if (sel) begin
      lineBuffer_5996 <= lineBuffer_5995;
    end
    if (sel) begin
      lineBuffer_5997 <= lineBuffer_5996;
    end
    if (sel) begin
      lineBuffer_5998 <= lineBuffer_5997;
    end
    if (sel) begin
      lineBuffer_5999 <= lineBuffer_5998;
    end
    if (sel) begin
      lineBuffer_6000 <= lineBuffer_5999;
    end
    if (sel) begin
      lineBuffer_6001 <= lineBuffer_6000;
    end
    if (sel) begin
      lineBuffer_6002 <= lineBuffer_6001;
    end
    if (sel) begin
      lineBuffer_6003 <= lineBuffer_6002;
    end
    if (sel) begin
      lineBuffer_6004 <= lineBuffer_6003;
    end
    if (sel) begin
      lineBuffer_6005 <= lineBuffer_6004;
    end
    if (sel) begin
      lineBuffer_6006 <= lineBuffer_6005;
    end
    if (sel) begin
      lineBuffer_6007 <= lineBuffer_6006;
    end
    if (sel) begin
      lineBuffer_6008 <= lineBuffer_6007;
    end
    if (sel) begin
      lineBuffer_6009 <= lineBuffer_6008;
    end
    if (sel) begin
      lineBuffer_6010 <= lineBuffer_6009;
    end
    if (sel) begin
      lineBuffer_6011 <= lineBuffer_6010;
    end
    if (sel) begin
      lineBuffer_6012 <= lineBuffer_6011;
    end
    if (sel) begin
      lineBuffer_6013 <= lineBuffer_6012;
    end
    if (sel) begin
      lineBuffer_6014 <= lineBuffer_6013;
    end
    if (sel) begin
      lineBuffer_6015 <= lineBuffer_6014;
    end
    if (sel) begin
      lineBuffer_6016 <= lineBuffer_6015;
    end
    if (sel) begin
      lineBuffer_6017 <= lineBuffer_6016;
    end
    if (sel) begin
      lineBuffer_6018 <= lineBuffer_6017;
    end
    if (sel) begin
      lineBuffer_6019 <= lineBuffer_6018;
    end
    if (sel) begin
      lineBuffer_6020 <= lineBuffer_6019;
    end
    if (sel) begin
      lineBuffer_6021 <= lineBuffer_6020;
    end
    if (sel) begin
      lineBuffer_6022 <= lineBuffer_6021;
    end
    if (sel) begin
      lineBuffer_6023 <= lineBuffer_6022;
    end
    if (sel) begin
      lineBuffer_6024 <= lineBuffer_6023;
    end
    if (sel) begin
      lineBuffer_6025 <= lineBuffer_6024;
    end
    if (sel) begin
      lineBuffer_6026 <= lineBuffer_6025;
    end
    if (sel) begin
      lineBuffer_6027 <= lineBuffer_6026;
    end
    if (sel) begin
      lineBuffer_6028 <= lineBuffer_6027;
    end
    if (sel) begin
      lineBuffer_6029 <= lineBuffer_6028;
    end
    if (sel) begin
      lineBuffer_6030 <= lineBuffer_6029;
    end
    if (sel) begin
      lineBuffer_6031 <= lineBuffer_6030;
    end
    if (sel) begin
      lineBuffer_6032 <= lineBuffer_6031;
    end
    if (sel) begin
      lineBuffer_6033 <= lineBuffer_6032;
    end
    if (sel) begin
      lineBuffer_6034 <= lineBuffer_6033;
    end
    if (sel) begin
      lineBuffer_6035 <= lineBuffer_6034;
    end
    if (sel) begin
      lineBuffer_6036 <= lineBuffer_6035;
    end
    if (sel) begin
      lineBuffer_6037 <= lineBuffer_6036;
    end
    if (sel) begin
      lineBuffer_6038 <= lineBuffer_6037;
    end
    if (sel) begin
      lineBuffer_6039 <= lineBuffer_6038;
    end
    if (sel) begin
      lineBuffer_6040 <= lineBuffer_6039;
    end
    if (sel) begin
      lineBuffer_6041 <= lineBuffer_6040;
    end
    if (sel) begin
      lineBuffer_6042 <= lineBuffer_6041;
    end
    if (sel) begin
      lineBuffer_6043 <= lineBuffer_6042;
    end
    if (sel) begin
      lineBuffer_6044 <= lineBuffer_6043;
    end
    if (sel) begin
      lineBuffer_6045 <= lineBuffer_6044;
    end
    if (sel) begin
      lineBuffer_6046 <= lineBuffer_6045;
    end
    if (sel) begin
      lineBuffer_6047 <= lineBuffer_6046;
    end
    if (sel) begin
      lineBuffer_6048 <= lineBuffer_6047;
    end
    if (sel) begin
      lineBuffer_6049 <= lineBuffer_6048;
    end
    if (sel) begin
      lineBuffer_6050 <= lineBuffer_6049;
    end
    if (sel) begin
      lineBuffer_6051 <= lineBuffer_6050;
    end
    if (sel) begin
      lineBuffer_6052 <= lineBuffer_6051;
    end
    if (sel) begin
      lineBuffer_6053 <= lineBuffer_6052;
    end
    if (sel) begin
      lineBuffer_6054 <= lineBuffer_6053;
    end
    if (sel) begin
      lineBuffer_6055 <= lineBuffer_6054;
    end
    if (sel) begin
      lineBuffer_6056 <= lineBuffer_6055;
    end
    if (sel) begin
      lineBuffer_6057 <= lineBuffer_6056;
    end
    if (sel) begin
      lineBuffer_6058 <= lineBuffer_6057;
    end
    if (sel) begin
      lineBuffer_6059 <= lineBuffer_6058;
    end
    if (sel) begin
      lineBuffer_6060 <= lineBuffer_6059;
    end
    if (sel) begin
      lineBuffer_6061 <= lineBuffer_6060;
    end
    if (sel) begin
      lineBuffer_6062 <= lineBuffer_6061;
    end
    if (sel) begin
      lineBuffer_6063 <= lineBuffer_6062;
    end
    if (sel) begin
      lineBuffer_6064 <= lineBuffer_6063;
    end
    if (sel) begin
      lineBuffer_6065 <= lineBuffer_6064;
    end
    if (sel) begin
      lineBuffer_6066 <= lineBuffer_6065;
    end
    if (sel) begin
      lineBuffer_6067 <= lineBuffer_6066;
    end
    if (sel) begin
      lineBuffer_6068 <= lineBuffer_6067;
    end
    if (sel) begin
      lineBuffer_6069 <= lineBuffer_6068;
    end
    if (sel) begin
      lineBuffer_6070 <= lineBuffer_6069;
    end
    if (sel) begin
      lineBuffer_6071 <= lineBuffer_6070;
    end
    if (sel) begin
      lineBuffer_6072 <= lineBuffer_6071;
    end
    if (sel) begin
      lineBuffer_6073 <= lineBuffer_6072;
    end
    if (sel) begin
      lineBuffer_6074 <= lineBuffer_6073;
    end
    if (sel) begin
      lineBuffer_6075 <= lineBuffer_6074;
    end
    if (sel) begin
      lineBuffer_6076 <= lineBuffer_6075;
    end
    if (sel) begin
      lineBuffer_6077 <= lineBuffer_6076;
    end
    if (sel) begin
      lineBuffer_6078 <= lineBuffer_6077;
    end
    if (sel) begin
      lineBuffer_6079 <= lineBuffer_6078;
    end
    if (sel) begin
      lineBuffer_6080 <= lineBuffer_6079;
    end
    if (sel) begin
      lineBuffer_6081 <= lineBuffer_6080;
    end
    if (sel) begin
      lineBuffer_6082 <= lineBuffer_6081;
    end
    if (sel) begin
      lineBuffer_6083 <= lineBuffer_6082;
    end
    if (sel) begin
      lineBuffer_6084 <= lineBuffer_6083;
    end
    if (sel) begin
      lineBuffer_6085 <= lineBuffer_6084;
    end
    if (sel) begin
      lineBuffer_6086 <= lineBuffer_6085;
    end
    if (sel) begin
      lineBuffer_6087 <= lineBuffer_6086;
    end
    if (sel) begin
      lineBuffer_6088 <= lineBuffer_6087;
    end
    if (sel) begin
      lineBuffer_6089 <= lineBuffer_6088;
    end
    if (sel) begin
      lineBuffer_6090 <= lineBuffer_6089;
    end
    if (sel) begin
      lineBuffer_6091 <= lineBuffer_6090;
    end
    if (sel) begin
      lineBuffer_6092 <= lineBuffer_6091;
    end
    if (sel) begin
      lineBuffer_6093 <= lineBuffer_6092;
    end
    if (sel) begin
      lineBuffer_6094 <= lineBuffer_6093;
    end
    if (sel) begin
      lineBuffer_6095 <= lineBuffer_6094;
    end
    if (sel) begin
      lineBuffer_6096 <= lineBuffer_6095;
    end
    if (sel) begin
      lineBuffer_6097 <= lineBuffer_6096;
    end
    if (sel) begin
      lineBuffer_6098 <= lineBuffer_6097;
    end
    if (sel) begin
      lineBuffer_6099 <= lineBuffer_6098;
    end
    if (sel) begin
      lineBuffer_6100 <= lineBuffer_6099;
    end
    if (sel) begin
      lineBuffer_6101 <= lineBuffer_6100;
    end
    if (sel) begin
      lineBuffer_6102 <= lineBuffer_6101;
    end
    if (sel) begin
      lineBuffer_6103 <= lineBuffer_6102;
    end
    if (sel) begin
      lineBuffer_6104 <= lineBuffer_6103;
    end
    if (sel) begin
      lineBuffer_6105 <= lineBuffer_6104;
    end
    if (sel) begin
      lineBuffer_6106 <= lineBuffer_6105;
    end
    if (sel) begin
      lineBuffer_6107 <= lineBuffer_6106;
    end
    if (sel) begin
      lineBuffer_6108 <= lineBuffer_6107;
    end
    if (sel) begin
      lineBuffer_6109 <= lineBuffer_6108;
    end
    if (sel) begin
      lineBuffer_6110 <= lineBuffer_6109;
    end
    if (sel) begin
      lineBuffer_6111 <= lineBuffer_6110;
    end
    if (sel) begin
      lineBuffer_6112 <= lineBuffer_6111;
    end
    if (sel) begin
      lineBuffer_6113 <= lineBuffer_6112;
    end
    if (sel) begin
      lineBuffer_6114 <= lineBuffer_6113;
    end
    if (sel) begin
      lineBuffer_6115 <= lineBuffer_6114;
    end
    if (sel) begin
      lineBuffer_6116 <= lineBuffer_6115;
    end
    if (sel) begin
      lineBuffer_6117 <= lineBuffer_6116;
    end
    if (sel) begin
      lineBuffer_6118 <= lineBuffer_6117;
    end
    if (sel) begin
      lineBuffer_6119 <= lineBuffer_6118;
    end
    if (sel) begin
      lineBuffer_6120 <= lineBuffer_6119;
    end
    if (sel) begin
      lineBuffer_6121 <= lineBuffer_6120;
    end
    if (sel) begin
      lineBuffer_6122 <= lineBuffer_6121;
    end
    if (sel) begin
      lineBuffer_6123 <= lineBuffer_6122;
    end
    if (sel) begin
      lineBuffer_6124 <= lineBuffer_6123;
    end
    if (sel) begin
      lineBuffer_6125 <= lineBuffer_6124;
    end
    if (sel) begin
      lineBuffer_6126 <= lineBuffer_6125;
    end
    if (sel) begin
      lineBuffer_6127 <= lineBuffer_6126;
    end
    if (sel) begin
      lineBuffer_6128 <= lineBuffer_6127;
    end
    if (sel) begin
      lineBuffer_6129 <= lineBuffer_6128;
    end
    if (sel) begin
      lineBuffer_6130 <= lineBuffer_6129;
    end
    if (sel) begin
      lineBuffer_6131 <= lineBuffer_6130;
    end
    if (sel) begin
      lineBuffer_6132 <= lineBuffer_6131;
    end
    if (sel) begin
      lineBuffer_6133 <= lineBuffer_6132;
    end
    if (sel) begin
      lineBuffer_6134 <= lineBuffer_6133;
    end
    if (sel) begin
      lineBuffer_6135 <= lineBuffer_6134;
    end
    if (sel) begin
      lineBuffer_6136 <= lineBuffer_6135;
    end
    if (sel) begin
      lineBuffer_6137 <= lineBuffer_6136;
    end
    if (sel) begin
      lineBuffer_6138 <= lineBuffer_6137;
    end
    if (sel) begin
      lineBuffer_6139 <= lineBuffer_6138;
    end
    if (sel) begin
      lineBuffer_6140 <= lineBuffer_6139;
    end
    if (sel) begin
      lineBuffer_6141 <= lineBuffer_6140;
    end
    if (sel) begin
      lineBuffer_6142 <= lineBuffer_6141;
    end
    if (sel) begin
      lineBuffer_6143 <= lineBuffer_6142;
    end
    if (sel) begin
      lineBuffer_6144 <= lineBuffer_6143;
    end
    if (sel) begin
      lineBuffer_6145 <= lineBuffer_6144;
    end
    if (sel) begin
      lineBuffer_6146 <= lineBuffer_6145;
    end
    if (sel) begin
      lineBuffer_6147 <= lineBuffer_6146;
    end
    if (sel) begin
      lineBuffer_6148 <= lineBuffer_6147;
    end
    if (sel) begin
      lineBuffer_6149 <= lineBuffer_6148;
    end
    if (sel) begin
      lineBuffer_6150 <= lineBuffer_6149;
    end
    if (sel) begin
      lineBuffer_6151 <= lineBuffer_6150;
    end
    if (sel) begin
      lineBuffer_6152 <= lineBuffer_6151;
    end
    if (sel) begin
      lineBuffer_6153 <= lineBuffer_6152;
    end
    if (sel) begin
      lineBuffer_6154 <= lineBuffer_6153;
    end
    if (sel) begin
      lineBuffer_6155 <= lineBuffer_6154;
    end
    if (sel) begin
      lineBuffer_6156 <= lineBuffer_6155;
    end
    if (sel) begin
      lineBuffer_6157 <= lineBuffer_6156;
    end
    if (sel) begin
      lineBuffer_6158 <= lineBuffer_6157;
    end
    if (sel) begin
      lineBuffer_6159 <= lineBuffer_6158;
    end
    if (sel) begin
      lineBuffer_6160 <= lineBuffer_6159;
    end
    if (sel) begin
      lineBuffer_6161 <= lineBuffer_6160;
    end
    if (sel) begin
      lineBuffer_6162 <= lineBuffer_6161;
    end
    if (sel) begin
      lineBuffer_6163 <= lineBuffer_6162;
    end
    if (sel) begin
      lineBuffer_6164 <= lineBuffer_6163;
    end
    if (sel) begin
      lineBuffer_6165 <= lineBuffer_6164;
    end
    if (sel) begin
      lineBuffer_6166 <= lineBuffer_6165;
    end
    if (sel) begin
      lineBuffer_6167 <= lineBuffer_6166;
    end
    if (sel) begin
      lineBuffer_6168 <= lineBuffer_6167;
    end
    if (sel) begin
      lineBuffer_6169 <= lineBuffer_6168;
    end
    if (sel) begin
      lineBuffer_6170 <= lineBuffer_6169;
    end
    if (sel) begin
      lineBuffer_6171 <= lineBuffer_6170;
    end
    if (sel) begin
      lineBuffer_6172 <= lineBuffer_6171;
    end
    if (sel) begin
      lineBuffer_6173 <= lineBuffer_6172;
    end
    if (sel) begin
      lineBuffer_6174 <= lineBuffer_6173;
    end
    if (sel) begin
      lineBuffer_6175 <= lineBuffer_6174;
    end
    if (sel) begin
      lineBuffer_6176 <= lineBuffer_6175;
    end
    if (sel) begin
      lineBuffer_6177 <= lineBuffer_6176;
    end
    if (sel) begin
      lineBuffer_6178 <= lineBuffer_6177;
    end
    if (sel) begin
      lineBuffer_6179 <= lineBuffer_6178;
    end
    if (sel) begin
      lineBuffer_6180 <= lineBuffer_6179;
    end
    if (sel) begin
      lineBuffer_6181 <= lineBuffer_6180;
    end
    if (sel) begin
      lineBuffer_6182 <= lineBuffer_6181;
    end
    if (sel) begin
      lineBuffer_6183 <= lineBuffer_6182;
    end
    if (sel) begin
      lineBuffer_6184 <= lineBuffer_6183;
    end
    if (sel) begin
      lineBuffer_6185 <= lineBuffer_6184;
    end
    if (sel) begin
      lineBuffer_6186 <= lineBuffer_6185;
    end
    if (sel) begin
      lineBuffer_6187 <= lineBuffer_6186;
    end
    if (sel) begin
      lineBuffer_6188 <= lineBuffer_6187;
    end
    if (sel) begin
      lineBuffer_6189 <= lineBuffer_6188;
    end
    if (sel) begin
      lineBuffer_6190 <= lineBuffer_6189;
    end
    if (sel) begin
      lineBuffer_6191 <= lineBuffer_6190;
    end
    if (sel) begin
      lineBuffer_6192 <= lineBuffer_6191;
    end
    if (sel) begin
      lineBuffer_6193 <= lineBuffer_6192;
    end
    if (sel) begin
      lineBuffer_6194 <= lineBuffer_6193;
    end
    if (sel) begin
      lineBuffer_6195 <= lineBuffer_6194;
    end
    if (sel) begin
      lineBuffer_6196 <= lineBuffer_6195;
    end
    if (sel) begin
      lineBuffer_6197 <= lineBuffer_6196;
    end
    if (sel) begin
      lineBuffer_6198 <= lineBuffer_6197;
    end
    if (sel) begin
      lineBuffer_6199 <= lineBuffer_6198;
    end
    if (sel) begin
      lineBuffer_6200 <= lineBuffer_6199;
    end
    if (sel) begin
      lineBuffer_6201 <= lineBuffer_6200;
    end
    if (sel) begin
      lineBuffer_6202 <= lineBuffer_6201;
    end
    if (sel) begin
      lineBuffer_6203 <= lineBuffer_6202;
    end
    if (sel) begin
      lineBuffer_6204 <= lineBuffer_6203;
    end
    if (sel) begin
      lineBuffer_6205 <= lineBuffer_6204;
    end
    if (sel) begin
      lineBuffer_6206 <= lineBuffer_6205;
    end
    if (sel) begin
      lineBuffer_6207 <= lineBuffer_6206;
    end
    if (sel) begin
      lineBuffer_6208 <= lineBuffer_6207;
    end
    if (sel) begin
      lineBuffer_6209 <= lineBuffer_6208;
    end
    if (sel) begin
      lineBuffer_6210 <= lineBuffer_6209;
    end
    if (sel) begin
      lineBuffer_6211 <= lineBuffer_6210;
    end
    if (sel) begin
      lineBuffer_6212 <= lineBuffer_6211;
    end
    if (sel) begin
      lineBuffer_6213 <= lineBuffer_6212;
    end
    if (sel) begin
      lineBuffer_6214 <= lineBuffer_6213;
    end
    if (sel) begin
      lineBuffer_6215 <= lineBuffer_6214;
    end
    if (sel) begin
      lineBuffer_6216 <= lineBuffer_6215;
    end
    if (sel) begin
      lineBuffer_6217 <= lineBuffer_6216;
    end
    if (sel) begin
      lineBuffer_6218 <= lineBuffer_6217;
    end
    if (sel) begin
      lineBuffer_6219 <= lineBuffer_6218;
    end
    if (sel) begin
      lineBuffer_6220 <= lineBuffer_6219;
    end
    if (sel) begin
      lineBuffer_6221 <= lineBuffer_6220;
    end
    if (sel) begin
      lineBuffer_6222 <= lineBuffer_6221;
    end
    if (sel) begin
      lineBuffer_6223 <= lineBuffer_6222;
    end
    if (sel) begin
      lineBuffer_6224 <= lineBuffer_6223;
    end
    if (sel) begin
      lineBuffer_6225 <= lineBuffer_6224;
    end
    if (sel) begin
      lineBuffer_6226 <= lineBuffer_6225;
    end
    if (sel) begin
      lineBuffer_6227 <= lineBuffer_6226;
    end
    if (sel) begin
      lineBuffer_6228 <= lineBuffer_6227;
    end
    if (sel) begin
      lineBuffer_6229 <= lineBuffer_6228;
    end
    if (sel) begin
      lineBuffer_6230 <= lineBuffer_6229;
    end
    if (sel) begin
      lineBuffer_6231 <= lineBuffer_6230;
    end
    if (sel) begin
      lineBuffer_6232 <= lineBuffer_6231;
    end
    if (sel) begin
      lineBuffer_6233 <= lineBuffer_6232;
    end
    if (sel) begin
      lineBuffer_6234 <= lineBuffer_6233;
    end
    if (sel) begin
      lineBuffer_6235 <= lineBuffer_6234;
    end
    if (sel) begin
      lineBuffer_6236 <= lineBuffer_6235;
    end
    if (sel) begin
      lineBuffer_6237 <= lineBuffer_6236;
    end
    if (sel) begin
      lineBuffer_6238 <= lineBuffer_6237;
    end
    if (sel) begin
      lineBuffer_6239 <= lineBuffer_6238;
    end
    if (sel) begin
      lineBuffer_6240 <= lineBuffer_6239;
    end
    if (sel) begin
      lineBuffer_6241 <= lineBuffer_6240;
    end
    if (sel) begin
      lineBuffer_6242 <= lineBuffer_6241;
    end
    if (sel) begin
      lineBuffer_6243 <= lineBuffer_6242;
    end
    if (sel) begin
      lineBuffer_6244 <= lineBuffer_6243;
    end
    if (sel) begin
      lineBuffer_6245 <= lineBuffer_6244;
    end
    if (sel) begin
      lineBuffer_6246 <= lineBuffer_6245;
    end
    if (sel) begin
      lineBuffer_6247 <= lineBuffer_6246;
    end
    if (sel) begin
      lineBuffer_6248 <= lineBuffer_6247;
    end
    if (sel) begin
      lineBuffer_6249 <= lineBuffer_6248;
    end
    if (sel) begin
      lineBuffer_6250 <= lineBuffer_6249;
    end
    if (sel) begin
      lineBuffer_6251 <= lineBuffer_6250;
    end
    if (sel) begin
      lineBuffer_6252 <= lineBuffer_6251;
    end
    if (sel) begin
      lineBuffer_6253 <= lineBuffer_6252;
    end
    if (sel) begin
      lineBuffer_6254 <= lineBuffer_6253;
    end
    if (sel) begin
      lineBuffer_6255 <= lineBuffer_6254;
    end
    if (sel) begin
      lineBuffer_6256 <= lineBuffer_6255;
    end
    if (sel) begin
      lineBuffer_6257 <= lineBuffer_6256;
    end
    if (sel) begin
      lineBuffer_6258 <= lineBuffer_6257;
    end
    if (sel) begin
      lineBuffer_6259 <= lineBuffer_6258;
    end
    if (sel) begin
      lineBuffer_6260 <= lineBuffer_6259;
    end
    if (sel) begin
      lineBuffer_6261 <= lineBuffer_6260;
    end
    if (sel) begin
      lineBuffer_6262 <= lineBuffer_6261;
    end
    if (sel) begin
      lineBuffer_6263 <= lineBuffer_6262;
    end
    if (sel) begin
      lineBuffer_6264 <= lineBuffer_6263;
    end
    if (sel) begin
      lineBuffer_6265 <= lineBuffer_6264;
    end
    if (sel) begin
      lineBuffer_6266 <= lineBuffer_6265;
    end
    if (sel) begin
      lineBuffer_6267 <= lineBuffer_6266;
    end
    if (sel) begin
      lineBuffer_6268 <= lineBuffer_6267;
    end
    if (sel) begin
      lineBuffer_6269 <= lineBuffer_6268;
    end
    if (sel) begin
      lineBuffer_6270 <= lineBuffer_6269;
    end
    if (sel) begin
      lineBuffer_6271 <= lineBuffer_6270;
    end
    if (sel) begin
      lineBuffer_6272 <= lineBuffer_6271;
    end
    if (sel) begin
      lineBuffer_6273 <= lineBuffer_6272;
    end
    if (sel) begin
      lineBuffer_6274 <= lineBuffer_6273;
    end
    if (sel) begin
      lineBuffer_6275 <= lineBuffer_6274;
    end
    if (sel) begin
      lineBuffer_6276 <= lineBuffer_6275;
    end
    if (sel) begin
      lineBuffer_6277 <= lineBuffer_6276;
    end
    if (sel) begin
      lineBuffer_6278 <= lineBuffer_6277;
    end
    if (sel) begin
      lineBuffer_6279 <= lineBuffer_6278;
    end
    if (sel) begin
      lineBuffer_6280 <= lineBuffer_6279;
    end
    if (sel) begin
      lineBuffer_6281 <= lineBuffer_6280;
    end
    if (sel) begin
      lineBuffer_6282 <= lineBuffer_6281;
    end
    if (sel) begin
      lineBuffer_6283 <= lineBuffer_6282;
    end
    if (sel) begin
      lineBuffer_6284 <= lineBuffer_6283;
    end
    if (sel) begin
      lineBuffer_6285 <= lineBuffer_6284;
    end
    if (sel) begin
      lineBuffer_6286 <= lineBuffer_6285;
    end
    if (sel) begin
      lineBuffer_6287 <= lineBuffer_6286;
    end
    if (sel) begin
      lineBuffer_6288 <= lineBuffer_6287;
    end
    if (sel) begin
      lineBuffer_6289 <= lineBuffer_6288;
    end
    if (sel) begin
      lineBuffer_6290 <= lineBuffer_6289;
    end
    if (sel) begin
      lineBuffer_6291 <= lineBuffer_6290;
    end
    if (sel) begin
      lineBuffer_6292 <= lineBuffer_6291;
    end
    if (sel) begin
      lineBuffer_6293 <= lineBuffer_6292;
    end
    if (sel) begin
      lineBuffer_6294 <= lineBuffer_6293;
    end
    if (sel) begin
      lineBuffer_6295 <= lineBuffer_6294;
    end
    if (sel) begin
      lineBuffer_6296 <= lineBuffer_6295;
    end
    if (sel) begin
      lineBuffer_6297 <= lineBuffer_6296;
    end
    if (sel) begin
      lineBuffer_6298 <= lineBuffer_6297;
    end
    if (sel) begin
      lineBuffer_6299 <= lineBuffer_6298;
    end
    if (sel) begin
      lineBuffer_6300 <= lineBuffer_6299;
    end
    if (sel) begin
      lineBuffer_6301 <= lineBuffer_6300;
    end
    if (sel) begin
      lineBuffer_6302 <= lineBuffer_6301;
    end
    if (sel) begin
      lineBuffer_6303 <= lineBuffer_6302;
    end
    if (sel) begin
      lineBuffer_6304 <= lineBuffer_6303;
    end
    if (sel) begin
      lineBuffer_6305 <= lineBuffer_6304;
    end
    if (sel) begin
      lineBuffer_6306 <= lineBuffer_6305;
    end
    if (sel) begin
      lineBuffer_6307 <= lineBuffer_6306;
    end
    if (sel) begin
      lineBuffer_6308 <= lineBuffer_6307;
    end
    if (sel) begin
      lineBuffer_6309 <= lineBuffer_6308;
    end
    if (sel) begin
      lineBuffer_6310 <= lineBuffer_6309;
    end
    if (sel) begin
      lineBuffer_6311 <= lineBuffer_6310;
    end
    if (sel) begin
      lineBuffer_6312 <= lineBuffer_6311;
    end
    if (sel) begin
      lineBuffer_6313 <= lineBuffer_6312;
    end
    if (sel) begin
      lineBuffer_6314 <= lineBuffer_6313;
    end
    if (sel) begin
      lineBuffer_6315 <= lineBuffer_6314;
    end
    if (sel) begin
      lineBuffer_6316 <= lineBuffer_6315;
    end
    if (sel) begin
      lineBuffer_6317 <= lineBuffer_6316;
    end
    if (sel) begin
      lineBuffer_6318 <= lineBuffer_6317;
    end
    if (sel) begin
      lineBuffer_6319 <= lineBuffer_6318;
    end
    if (sel) begin
      lineBuffer_6320 <= lineBuffer_6319;
    end
    if (sel) begin
      lineBuffer_6321 <= lineBuffer_6320;
    end
    if (sel) begin
      lineBuffer_6322 <= lineBuffer_6321;
    end
    if (sel) begin
      lineBuffer_6323 <= lineBuffer_6322;
    end
    if (sel) begin
      lineBuffer_6324 <= lineBuffer_6323;
    end
    if (sel) begin
      lineBuffer_6325 <= lineBuffer_6324;
    end
    if (sel) begin
      lineBuffer_6326 <= lineBuffer_6325;
    end
    if (sel) begin
      lineBuffer_6327 <= lineBuffer_6326;
    end
    if (sel) begin
      lineBuffer_6328 <= lineBuffer_6327;
    end
    if (sel) begin
      lineBuffer_6329 <= lineBuffer_6328;
    end
    if (sel) begin
      lineBuffer_6330 <= lineBuffer_6329;
    end
    if (sel) begin
      lineBuffer_6331 <= lineBuffer_6330;
    end
    if (sel) begin
      lineBuffer_6332 <= lineBuffer_6331;
    end
    if (sel) begin
      lineBuffer_6333 <= lineBuffer_6332;
    end
    if (sel) begin
      lineBuffer_6334 <= lineBuffer_6333;
    end
    if (sel) begin
      lineBuffer_6335 <= lineBuffer_6334;
    end
    if (sel) begin
      lineBuffer_6336 <= lineBuffer_6335;
    end
    if (sel) begin
      lineBuffer_6337 <= lineBuffer_6336;
    end
    if (sel) begin
      lineBuffer_6338 <= lineBuffer_6337;
    end
    if (sel) begin
      lineBuffer_6339 <= lineBuffer_6338;
    end
    if (sel) begin
      lineBuffer_6340 <= lineBuffer_6339;
    end
    if (sel) begin
      lineBuffer_6341 <= lineBuffer_6340;
    end
    if (sel) begin
      lineBuffer_6342 <= lineBuffer_6341;
    end
    if (sel) begin
      lineBuffer_6343 <= lineBuffer_6342;
    end
    if (sel) begin
      lineBuffer_6344 <= lineBuffer_6343;
    end
    if (sel) begin
      lineBuffer_6345 <= lineBuffer_6344;
    end
    if (sel) begin
      lineBuffer_6346 <= lineBuffer_6345;
    end
    if (sel) begin
      lineBuffer_6347 <= lineBuffer_6346;
    end
    if (sel) begin
      lineBuffer_6348 <= lineBuffer_6347;
    end
    if (sel) begin
      lineBuffer_6349 <= lineBuffer_6348;
    end
    if (sel) begin
      lineBuffer_6350 <= lineBuffer_6349;
    end
    if (sel) begin
      lineBuffer_6351 <= lineBuffer_6350;
    end
    if (sel) begin
      lineBuffer_6352 <= lineBuffer_6351;
    end
    if (sel) begin
      lineBuffer_6353 <= lineBuffer_6352;
    end
    if (sel) begin
      lineBuffer_6354 <= lineBuffer_6353;
    end
    if (sel) begin
      lineBuffer_6355 <= lineBuffer_6354;
    end
    if (sel) begin
      lineBuffer_6356 <= lineBuffer_6355;
    end
    if (sel) begin
      lineBuffer_6357 <= lineBuffer_6356;
    end
    if (sel) begin
      lineBuffer_6358 <= lineBuffer_6357;
    end
    if (sel) begin
      lineBuffer_6359 <= lineBuffer_6358;
    end
    if (sel) begin
      lineBuffer_6360 <= lineBuffer_6359;
    end
    if (sel) begin
      lineBuffer_6361 <= lineBuffer_6360;
    end
    if (sel) begin
      lineBuffer_6362 <= lineBuffer_6361;
    end
    if (sel) begin
      lineBuffer_6363 <= lineBuffer_6362;
    end
    if (sel) begin
      lineBuffer_6364 <= lineBuffer_6363;
    end
    if (sel) begin
      lineBuffer_6365 <= lineBuffer_6364;
    end
    if (sel) begin
      lineBuffer_6366 <= lineBuffer_6365;
    end
    if (sel) begin
      lineBuffer_6367 <= lineBuffer_6366;
    end
    if (sel) begin
      lineBuffer_6368 <= lineBuffer_6367;
    end
    if (sel) begin
      lineBuffer_6369 <= lineBuffer_6368;
    end
    if (sel) begin
      lineBuffer_6370 <= lineBuffer_6369;
    end
    if (sel) begin
      lineBuffer_6371 <= lineBuffer_6370;
    end
    if (sel) begin
      lineBuffer_6372 <= lineBuffer_6371;
    end
    if (sel) begin
      lineBuffer_6373 <= lineBuffer_6372;
    end
    if (sel) begin
      lineBuffer_6374 <= lineBuffer_6373;
    end
    if (sel) begin
      lineBuffer_6375 <= lineBuffer_6374;
    end
    if (sel) begin
      lineBuffer_6376 <= lineBuffer_6375;
    end
    if (sel) begin
      lineBuffer_6377 <= lineBuffer_6376;
    end
    if (sel) begin
      lineBuffer_6378 <= lineBuffer_6377;
    end
    if (sel) begin
      lineBuffer_6379 <= lineBuffer_6378;
    end
    if (sel) begin
      lineBuffer_6380 <= lineBuffer_6379;
    end
    if (sel) begin
      lineBuffer_6381 <= lineBuffer_6380;
    end
    if (sel) begin
      lineBuffer_6382 <= lineBuffer_6381;
    end
    if (sel) begin
      lineBuffer_6383 <= lineBuffer_6382;
    end
    if (sel) begin
      lineBuffer_6384 <= lineBuffer_6383;
    end
    if (sel) begin
      lineBuffer_6385 <= lineBuffer_6384;
    end
    if (sel) begin
      lineBuffer_6386 <= lineBuffer_6385;
    end
    if (sel) begin
      lineBuffer_6387 <= lineBuffer_6386;
    end
    if (sel) begin
      lineBuffer_6388 <= lineBuffer_6387;
    end
    if (sel) begin
      lineBuffer_6389 <= lineBuffer_6388;
    end
    if (sel) begin
      lineBuffer_6390 <= lineBuffer_6389;
    end
    if (sel) begin
      lineBuffer_6391 <= lineBuffer_6390;
    end
    if (sel) begin
      lineBuffer_6392 <= lineBuffer_6391;
    end
    if (sel) begin
      lineBuffer_6393 <= lineBuffer_6392;
    end
    if (sel) begin
      lineBuffer_6394 <= lineBuffer_6393;
    end
    if (sel) begin
      lineBuffer_6395 <= lineBuffer_6394;
    end
    if (sel) begin
      lineBuffer_6396 <= lineBuffer_6395;
    end
    if (sel) begin
      lineBuffer_6397 <= lineBuffer_6396;
    end
    if (sel) begin
      lineBuffer_6398 <= lineBuffer_6397;
    end
    if (sel) begin
      lineBuffer_6399 <= lineBuffer_6398;
    end
    if (sel) begin
      windowBuffer_0 <= windowBuffer_1;
    end
    if (sel) begin
      windowBuffer_1 <= windowBuffer_2;
    end
    if (sel) begin
      windowBuffer_2 <= windowBuffer_3;
    end
    if (sel) begin
      windowBuffer_3 <= windowBuffer_4;
    end
    if (sel) begin
      windowBuffer_4 <= lineBuffer_1279;
    end
    if (sel) begin
      windowBuffer_5 <= windowBuffer_6;
    end
    if (sel) begin
      windowBuffer_6 <= windowBuffer_7;
    end
    if (sel) begin
      windowBuffer_7 <= windowBuffer_8;
    end
    if (sel) begin
      windowBuffer_8 <= windowBuffer_9;
    end
    if (sel) begin
      windowBuffer_9 <= lineBuffer_2559;
    end
    if (sel) begin
      windowBuffer_10 <= windowBuffer_11;
    end
    if (sel) begin
      windowBuffer_11 <= windowBuffer_12;
    end
    if (sel) begin
      windowBuffer_12 <= windowBuffer_13;
    end
    if (sel) begin
      windowBuffer_13 <= windowBuffer_14;
    end
    if (sel) begin
      windowBuffer_14 <= lineBuffer_3839;
    end
    if (sel) begin
      windowBuffer_15 <= windowBuffer_16;
    end
    if (sel) begin
      windowBuffer_16 <= windowBuffer_17;
    end
    if (sel) begin
      windowBuffer_17 <= windowBuffer_18;
    end
    if (sel) begin
      windowBuffer_18 <= windowBuffer_19;
    end
    if (sel) begin
      windowBuffer_19 <= lineBuffer_5119;
    end
    if (sel) begin
      windowBuffer_20 <= windowBuffer_21;
    end
    if (sel) begin
      windowBuffer_21 <= windowBuffer_22;
    end
    if (sel) begin
      windowBuffer_22 <= windowBuffer_23;
    end
    if (sel) begin
      windowBuffer_23 <= windowBuffer_24;
    end
    if (sel) begin
      windowBuffer_24 <= lineBuffer_6399;
    end
  end
endmodule
module NothingFilter(
  input        clock,
  input        reset,
  output       io_enq_ready,
  input        io_enq_valid,
  input  [7:0] io_enq_bits,
  input        io_enq_user,
  input        io_enq_last,
  input        io_deq_ready,
  output       io_deq_valid,
  output [7:0] io_deq_bits,
  output       io_deq_user,
  output       io_deq_last
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
`endif // RANDOMIZE_REG_INIT
  reg [1:0] stateReg; // @[ChiselImProc.scala 56:28]
  reg [7:0] dataReg; // @[ChiselImProc.scala 58:23]
  reg [7:0] shadowReg; // @[ChiselImProc.scala 60:25]
  reg  userReg; // @[ChiselImProc.scala 61:23]
  reg  shadowUserReg; // @[ChiselImProc.scala 62:29]
  reg  lastReg; // @[ChiselImProc.scala 63:23]
  reg  shadowLastReg; // @[ChiselImProc.scala 64:29]
  wire  _T = 2'h0 == stateReg; // @[Conditional.scala 37:30]
  wire  _T_1 = 2'h1 == stateReg; // @[Conditional.scala 37:30]
  wire  _T_2 = ~io_enq_valid; // @[ChiselImProc.scala 78:39]
  wire  _T_3 = io_deq_ready & _T_2; // @[ChiselImProc.scala 78:36]
  wire  _T_4 = io_deq_ready & io_enq_valid; // @[ChiselImProc.scala 81:42]
  wire  _T_5 = ~io_deq_ready; // @[ChiselImProc.scala 86:29]
  wire  _T_6 = _T_5 & io_enq_valid; // @[ChiselImProc.scala 86:43]
  wire  _T_7 = 2'h2 == stateReg; // @[Conditional.scala 37:30]
  wire  _T_8 = 2'h3 == stateReg; // @[Conditional.scala 37:30]
  wire  _T_9 = stateReg == 2'h0; // @[ChiselImProc.scala 110:35]
  wire  _T_10 = stateReg == 2'h1; // @[ChiselImProc.scala 110:57]
  wire  _T_11 = _T_9 | _T_10; // @[ChiselImProc.scala 110:45]
  wire  _T_12 = stateReg == 2'h3; // @[ChiselImProc.scala 110:77]
  wire  _T_15 = stateReg == 2'h2; // @[ChiselImProc.scala 111:55]
  assign io_enq_ready = _T_11 | _T_12; // @[ChiselImProc.scala 110:22]
  assign io_deq_valid = _T_10 | _T_15; // @[ChiselImProc.scala 111:22]
  assign io_deq_bits = dataReg; // @[ChiselImProc.scala 146:17]
  assign io_deq_user = userReg; // @[ChiselImProc.scala 138:17 ChiselImProc.scala 108:21]
  assign io_deq_last = lastReg; // @[ChiselImProc.scala 137:17 ChiselImProc.scala 107:21]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  stateReg = _RAND_0[1:0];
  _RAND_1 = {1{`RANDOM}};
  dataReg = _RAND_1[7:0];
  _RAND_2 = {1{`RANDOM}};
  shadowReg = _RAND_2[7:0];
  _RAND_3 = {1{`RANDOM}};
  userReg = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  shadowUserReg = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  lastReg = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  shadowLastReg = _RAND_6[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      stateReg <= 2'h0;
    end else if (_T) begin
      if (io_enq_valid) begin
        stateReg <= 2'h1;
      end
    end else if (_T_1) begin
      if (_T_3) begin
        stateReg <= 2'h0;
      end else if (_T_4) begin
        stateReg <= 2'h1;
      end else if (_T_6) begin
        stateReg <= 2'h2;
      end
    end else if (_T_7) begin
      if (io_deq_ready) begin
        stateReg <= 2'h1;
      end
    end else if (_T_8) begin
      stateReg <= 2'h0;
    end
    if (_T) begin
      if (io_enq_valid) begin
        dataReg <= io_enq_bits;
      end
    end else if (_T_1) begin
      if (!(_T_3)) begin
        if (_T_4) begin
          dataReg <= io_enq_bits;
        end
      end
    end else if (_T_7) begin
      if (io_deq_ready) begin
        dataReg <= shadowReg;
      end
    end
    if (!(_T)) begin
      if (_T_1) begin
        if (!(_T_3)) begin
          if (!(_T_4)) begin
            if (_T_6) begin
              shadowReg <= io_enq_bits;
            end
          end
        end
      end
    end
    if (_T) begin
      userReg <= io_enq_user;
    end else if (_T_1) begin
      if (_T_3) begin
        userReg <= io_enq_user;
      end else if (_T_4) begin
        userReg <= io_enq_user;
      end
    end else if (_T_7) begin
      if (io_deq_ready) begin
        userReg <= shadowUserReg;
      end
    end
    if (!(_T)) begin
      if (_T_1) begin
        if (!(_T_3)) begin
          if (!(_T_4)) begin
            if (_T_6) begin
              shadowUserReg <= io_enq_user;
            end
          end
        end
      end
    end
    if (_T) begin
      if (io_enq_valid) begin
        lastReg <= io_enq_last;
      end
    end else if (_T_1) begin
      if (!(_T_3)) begin
        if (_T_4) begin
          lastReg <= io_enq_last;
        end
      end
    end else if (_T_7) begin
      if (io_deq_ready) begin
        lastReg <= shadowLastReg;
      end
    end
    if (!(_T)) begin
      if (_T_1) begin
        if (!(_T_3)) begin
          if (!(_T_4)) begin
            if (_T_6) begin
              shadowLastReg <= io_enq_last;
            end
          end
        end
      end
    end
  end
endmodule
module Gray2RGBFilter(
  input         clock,
  input         reset,
  output        io_enq_ready,
  input         io_enq_valid,
  input  [23:0] io_enq_bits,
  input         io_enq_user,
  input         io_enq_last,
  input         io_deq_ready,
  output        io_deq_valid,
  output [23:0] io_deq_bits,
  output        io_deq_user,
  output        io_deq_last
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
`endif // RANDOMIZE_REG_INIT
  reg [1:0] stateReg; // @[ChiselImProc.scala 56:28]
  reg [23:0] dataReg; // @[ChiselImProc.scala 58:23]
  reg [23:0] shadowReg; // @[ChiselImProc.scala 60:25]
  reg  userReg; // @[ChiselImProc.scala 61:23]
  reg  shadowUserReg; // @[ChiselImProc.scala 62:29]
  reg  lastReg; // @[ChiselImProc.scala 63:23]
  reg  shadowLastReg; // @[ChiselImProc.scala 64:29]
  wire  _T = 2'h0 == stateReg; // @[Conditional.scala 37:30]
  wire  _T_1 = 2'h1 == stateReg; // @[Conditional.scala 37:30]
  wire  _T_2 = ~io_enq_valid; // @[ChiselImProc.scala 78:39]
  wire  _T_3 = io_deq_ready & _T_2; // @[ChiselImProc.scala 78:36]
  wire  _T_4 = io_deq_ready & io_enq_valid; // @[ChiselImProc.scala 81:42]
  wire  _T_5 = ~io_deq_ready; // @[ChiselImProc.scala 86:29]
  wire  _T_6 = _T_5 & io_enq_valid; // @[ChiselImProc.scala 86:43]
  wire  _T_7 = 2'h2 == stateReg; // @[Conditional.scala 37:30]
  wire  _T_8 = 2'h3 == stateReg; // @[Conditional.scala 37:30]
  wire  _T_9 = stateReg == 2'h0; // @[ChiselImProc.scala 110:35]
  wire  _T_10 = stateReg == 2'h1; // @[ChiselImProc.scala 110:57]
  wire  _T_11 = _T_9 | _T_10; // @[ChiselImProc.scala 110:45]
  wire  _T_12 = stateReg == 2'h3; // @[ChiselImProc.scala 110:77]
  wire  _T_15 = stateReg == 2'h2; // @[ChiselImProc.scala 111:55]
  wire [39:0] _GEN_44 = {dataReg, 16'h0}; // @[ChiselImProc.scala 174:28]
  wire [54:0] _T_17 = {{15'd0}, _GEN_44}; // @[ChiselImProc.scala 174:28]
  wire [31:0] _GEN_45 = {dataReg, 8'h0}; // @[ChiselImProc.scala 174:46]
  wire [38:0] _T_18 = {{7'd0}, _GEN_45}; // @[ChiselImProc.scala 174:46]
  wire [54:0] _GEN_46 = {{16'd0}, _T_18}; // @[ChiselImProc.scala 174:36]
  wire [54:0] _T_19 = _T_17 | _GEN_46; // @[ChiselImProc.scala 174:36]
  wire [54:0] _GEN_47 = {{31'd0}, dataReg}; // @[ChiselImProc.scala 174:53]
  wire [54:0] _T_20 = _T_19 | _GEN_47; // @[ChiselImProc.scala 174:53]
  assign io_enq_ready = _T_11 | _T_12; // @[ChiselImProc.scala 110:22]
  assign io_deq_valid = _T_10 | _T_15; // @[ChiselImProc.scala 111:22]
  assign io_deq_bits = _T_20[23:0]; // @[ChiselImProc.scala 174:17]
  assign io_deq_user = userReg; // @[ChiselImProc.scala 138:17 ChiselImProc.scala 108:21]
  assign io_deq_last = lastReg; // @[ChiselImProc.scala 137:17 ChiselImProc.scala 107:21]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  stateReg = _RAND_0[1:0];
  _RAND_1 = {1{`RANDOM}};
  dataReg = _RAND_1[23:0];
  _RAND_2 = {1{`RANDOM}};
  shadowReg = _RAND_2[23:0];
  _RAND_3 = {1{`RANDOM}};
  userReg = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  shadowUserReg = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  lastReg = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  shadowLastReg = _RAND_6[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      stateReg <= 2'h0;
    end else if (_T) begin
      if (io_enq_valid) begin
        stateReg <= 2'h1;
      end
    end else if (_T_1) begin
      if (_T_3) begin
        stateReg <= 2'h0;
      end else if (_T_4) begin
        stateReg <= 2'h1;
      end else if (_T_6) begin
        stateReg <= 2'h2;
      end
    end else if (_T_7) begin
      if (io_deq_ready) begin
        stateReg <= 2'h1;
      end
    end else if (_T_8) begin
      stateReg <= 2'h0;
    end
    if (_T) begin
      if (io_enq_valid) begin
        dataReg <= io_enq_bits;
      end
    end else if (_T_1) begin
      if (!(_T_3)) begin
        if (_T_4) begin
          dataReg <= io_enq_bits;
        end
      end
    end else if (_T_7) begin
      if (io_deq_ready) begin
        dataReg <= shadowReg;
      end
    end
    if (!(_T)) begin
      if (_T_1) begin
        if (!(_T_3)) begin
          if (!(_T_4)) begin
            if (_T_6) begin
              shadowReg <= io_enq_bits;
            end
          end
        end
      end
    end
    if (_T) begin
      userReg <= io_enq_user;
    end else if (_T_1) begin
      if (_T_3) begin
        userReg <= io_enq_user;
      end else if (_T_4) begin
        userReg <= io_enq_user;
      end
    end else if (_T_7) begin
      if (io_deq_ready) begin
        userReg <= shadowUserReg;
      end
    end
    if (!(_T)) begin
      if (_T_1) begin
        if (!(_T_3)) begin
          if (!(_T_4)) begin
            if (_T_6) begin
              shadowUserReg <= io_enq_user;
            end
          end
        end
      end
    end
    if (_T) begin
      if (io_enq_valid) begin
        lastReg <= io_enq_last;
      end
    end else if (_T_1) begin
      if (!(_T_3)) begin
        if (_T_4) begin
          lastReg <= io_enq_last;
        end
      end
    end else if (_T_7) begin
      if (io_deq_ready) begin
        lastReg <= shadowLastReg;
      end
    end
    if (!(_T)) begin
      if (_T_1) begin
        if (!(_T_3)) begin
          if (!(_T_4)) begin
            if (_T_6) begin
              shadowLastReg <= io_enq_last;
            end
          end
        end
      end
    end
  end
endmodule
module ChiselImProc(
  input         clock,
  input         reset,
  output        io_enq_ready,
  input         io_enq_valid,
  input  [23:0] io_enq_bits,
  input         io_enq_user,
  input         io_enq_last,
  input         io_deq_ready,
  output        io_deq_valid,
  output [23:0] io_deq_bits,
  output        io_deq_user,
  output        io_deq_last,
  output [31:0] io_dport,
  output [31:0] io_dport2
);
  wire  RGB2GrayFilter_clock; // @[ChiselImProc.scala 456:16]
  wire  RGB2GrayFilter_reset; // @[ChiselImProc.scala 456:16]
  wire  RGB2GrayFilter_io_enq_ready; // @[ChiselImProc.scala 456:16]
  wire  RGB2GrayFilter_io_enq_valid; // @[ChiselImProc.scala 456:16]
  wire [23:0] RGB2GrayFilter_io_enq_bits; // @[ChiselImProc.scala 456:16]
  wire  RGB2GrayFilter_io_enq_user; // @[ChiselImProc.scala 456:16]
  wire  RGB2GrayFilter_io_enq_last; // @[ChiselImProc.scala 456:16]
  wire  RGB2GrayFilter_io_deq_ready; // @[ChiselImProc.scala 456:16]
  wire  RGB2GrayFilter_io_deq_valid; // @[ChiselImProc.scala 456:16]
  wire [23:0] RGB2GrayFilter_io_deq_bits; // @[ChiselImProc.scala 456:16]
  wire  RGB2GrayFilter_io_deq_user; // @[ChiselImProc.scala 456:16]
  wire  RGB2GrayFilter_io_deq_last; // @[ChiselImProc.scala 456:16]
  wire  GaussianBlurFilter_clock; // @[ChiselImProc.scala 458:16]
  wire  GaussianBlurFilter_reset; // @[ChiselImProc.scala 458:16]
  wire  GaussianBlurFilter_io_enq_ready; // @[ChiselImProc.scala 458:16]
  wire  GaussianBlurFilter_io_enq_valid; // @[ChiselImProc.scala 458:16]
  wire [7:0] GaussianBlurFilter_io_enq_bits; // @[ChiselImProc.scala 458:16]
  wire  GaussianBlurFilter_io_enq_user; // @[ChiselImProc.scala 458:16]
  wire  GaussianBlurFilter_io_enq_last; // @[ChiselImProc.scala 458:16]
  wire  GaussianBlurFilter_io_deq_ready; // @[ChiselImProc.scala 458:16]
  wire  GaussianBlurFilter_io_deq_valid; // @[ChiselImProc.scala 458:16]
  wire [7:0] GaussianBlurFilter_io_deq_bits; // @[ChiselImProc.scala 458:16]
  wire  GaussianBlurFilter_io_deq_user; // @[ChiselImProc.scala 458:16]
  wire  GaussianBlurFilter_io_deq_last; // @[ChiselImProc.scala 458:16]
  wire  NothingFilter_clock; // @[ChiselImProc.scala 462:16]
  wire  NothingFilter_reset; // @[ChiselImProc.scala 462:16]
  wire  NothingFilter_io_enq_ready; // @[ChiselImProc.scala 462:16]
  wire  NothingFilter_io_enq_valid; // @[ChiselImProc.scala 462:16]
  wire [7:0] NothingFilter_io_enq_bits; // @[ChiselImProc.scala 462:16]
  wire  NothingFilter_io_enq_user; // @[ChiselImProc.scala 462:16]
  wire  NothingFilter_io_enq_last; // @[ChiselImProc.scala 462:16]
  wire  NothingFilter_io_deq_ready; // @[ChiselImProc.scala 462:16]
  wire  NothingFilter_io_deq_valid; // @[ChiselImProc.scala 462:16]
  wire [7:0] NothingFilter_io_deq_bits; // @[ChiselImProc.scala 462:16]
  wire  NothingFilter_io_deq_user; // @[ChiselImProc.scala 462:16]
  wire  NothingFilter_io_deq_last; // @[ChiselImProc.scala 462:16]
  wire  NothingFilter_1_clock; // @[ChiselImProc.scala 466:16]
  wire  NothingFilter_1_reset; // @[ChiselImProc.scala 466:16]
  wire  NothingFilter_1_io_enq_ready; // @[ChiselImProc.scala 466:16]
  wire  NothingFilter_1_io_enq_valid; // @[ChiselImProc.scala 466:16]
  wire [7:0] NothingFilter_1_io_enq_bits; // @[ChiselImProc.scala 466:16]
  wire  NothingFilter_1_io_enq_user; // @[ChiselImProc.scala 466:16]
  wire  NothingFilter_1_io_enq_last; // @[ChiselImProc.scala 466:16]
  wire  NothingFilter_1_io_deq_ready; // @[ChiselImProc.scala 466:16]
  wire  NothingFilter_1_io_deq_valid; // @[ChiselImProc.scala 466:16]
  wire [7:0] NothingFilter_1_io_deq_bits; // @[ChiselImProc.scala 466:16]
  wire  NothingFilter_1_io_deq_user; // @[ChiselImProc.scala 466:16]
  wire  NothingFilter_1_io_deq_last; // @[ChiselImProc.scala 466:16]
  wire  NothingFilter_2_clock; // @[ChiselImProc.scala 469:16]
  wire  NothingFilter_2_reset; // @[ChiselImProc.scala 469:16]
  wire  NothingFilter_2_io_enq_ready; // @[ChiselImProc.scala 469:16]
  wire  NothingFilter_2_io_enq_valid; // @[ChiselImProc.scala 469:16]
  wire [7:0] NothingFilter_2_io_enq_bits; // @[ChiselImProc.scala 469:16]
  wire  NothingFilter_2_io_enq_user; // @[ChiselImProc.scala 469:16]
  wire  NothingFilter_2_io_enq_last; // @[ChiselImProc.scala 469:16]
  wire  NothingFilter_2_io_deq_ready; // @[ChiselImProc.scala 469:16]
  wire  NothingFilter_2_io_deq_valid; // @[ChiselImProc.scala 469:16]
  wire [7:0] NothingFilter_2_io_deq_bits; // @[ChiselImProc.scala 469:16]
  wire  NothingFilter_2_io_deq_user; // @[ChiselImProc.scala 469:16]
  wire  NothingFilter_2_io_deq_last; // @[ChiselImProc.scala 469:16]
  wire  NothingFilter_3_clock; // @[ChiselImProc.scala 472:16]
  wire  NothingFilter_3_reset; // @[ChiselImProc.scala 472:16]
  wire  NothingFilter_3_io_enq_ready; // @[ChiselImProc.scala 472:16]
  wire  NothingFilter_3_io_enq_valid; // @[ChiselImProc.scala 472:16]
  wire [7:0] NothingFilter_3_io_enq_bits; // @[ChiselImProc.scala 472:16]
  wire  NothingFilter_3_io_enq_user; // @[ChiselImProc.scala 472:16]
  wire  NothingFilter_3_io_enq_last; // @[ChiselImProc.scala 472:16]
  wire  NothingFilter_3_io_deq_ready; // @[ChiselImProc.scala 472:16]
  wire  NothingFilter_3_io_deq_valid; // @[ChiselImProc.scala 472:16]
  wire [7:0] NothingFilter_3_io_deq_bits; // @[ChiselImProc.scala 472:16]
  wire  NothingFilter_3_io_deq_user; // @[ChiselImProc.scala 472:16]
  wire  NothingFilter_3_io_deq_last; // @[ChiselImProc.scala 472:16]
  wire  Gray2RGBFilter_clock; // @[ChiselImProc.scala 474:16]
  wire  Gray2RGBFilter_reset; // @[ChiselImProc.scala 474:16]
  wire  Gray2RGBFilter_io_enq_ready; // @[ChiselImProc.scala 474:16]
  wire  Gray2RGBFilter_io_enq_valid; // @[ChiselImProc.scala 474:16]
  wire [23:0] Gray2RGBFilter_io_enq_bits; // @[ChiselImProc.scala 474:16]
  wire  Gray2RGBFilter_io_enq_user; // @[ChiselImProc.scala 474:16]
  wire  Gray2RGBFilter_io_enq_last; // @[ChiselImProc.scala 474:16]
  wire  Gray2RGBFilter_io_deq_ready; // @[ChiselImProc.scala 474:16]
  wire  Gray2RGBFilter_io_deq_valid; // @[ChiselImProc.scala 474:16]
  wire [23:0] Gray2RGBFilter_io_deq_bits; // @[ChiselImProc.scala 474:16]
  wire  Gray2RGBFilter_io_deq_user; // @[ChiselImProc.scala 474:16]
  wire  Gray2RGBFilter_io_deq_last; // @[ChiselImProc.scala 474:16]
  RGB2GrayFilter RGB2GrayFilter ( // @[ChiselImProc.scala 456:16]
    .clock(RGB2GrayFilter_clock),
    .reset(RGB2GrayFilter_reset),
    .io_enq_ready(RGB2GrayFilter_io_enq_ready),
    .io_enq_valid(RGB2GrayFilter_io_enq_valid),
    .io_enq_bits(RGB2GrayFilter_io_enq_bits),
    .io_enq_user(RGB2GrayFilter_io_enq_user),
    .io_enq_last(RGB2GrayFilter_io_enq_last),
    .io_deq_ready(RGB2GrayFilter_io_deq_ready),
    .io_deq_valid(RGB2GrayFilter_io_deq_valid),
    .io_deq_bits(RGB2GrayFilter_io_deq_bits),
    .io_deq_user(RGB2GrayFilter_io_deq_user),
    .io_deq_last(RGB2GrayFilter_io_deq_last)
  );
  GaussianBlurFilter GaussianBlurFilter ( // @[ChiselImProc.scala 458:16]
    .clock(GaussianBlurFilter_clock),
    .reset(GaussianBlurFilter_reset),
    .io_enq_ready(GaussianBlurFilter_io_enq_ready),
    .io_enq_valid(GaussianBlurFilter_io_enq_valid),
    .io_enq_bits(GaussianBlurFilter_io_enq_bits),
    .io_enq_user(GaussianBlurFilter_io_enq_user),
    .io_enq_last(GaussianBlurFilter_io_enq_last),
    .io_deq_ready(GaussianBlurFilter_io_deq_ready),
    .io_deq_valid(GaussianBlurFilter_io_deq_valid),
    .io_deq_bits(GaussianBlurFilter_io_deq_bits),
    .io_deq_user(GaussianBlurFilter_io_deq_user),
    .io_deq_last(GaussianBlurFilter_io_deq_last)
  );
  NothingFilter NothingFilter ( // @[ChiselImProc.scala 462:16]
    .clock(NothingFilter_clock),
    .reset(NothingFilter_reset),
    .io_enq_ready(NothingFilter_io_enq_ready),
    .io_enq_valid(NothingFilter_io_enq_valid),
    .io_enq_bits(NothingFilter_io_enq_bits),
    .io_enq_user(NothingFilter_io_enq_user),
    .io_enq_last(NothingFilter_io_enq_last),
    .io_deq_ready(NothingFilter_io_deq_ready),
    .io_deq_valid(NothingFilter_io_deq_valid),
    .io_deq_bits(NothingFilter_io_deq_bits),
    .io_deq_user(NothingFilter_io_deq_user),
    .io_deq_last(NothingFilter_io_deq_last)
  );
  NothingFilter NothingFilter_1 ( // @[ChiselImProc.scala 466:16]
    .clock(NothingFilter_1_clock),
    .reset(NothingFilter_1_reset),
    .io_enq_ready(NothingFilter_1_io_enq_ready),
    .io_enq_valid(NothingFilter_1_io_enq_valid),
    .io_enq_bits(NothingFilter_1_io_enq_bits),
    .io_enq_user(NothingFilter_1_io_enq_user),
    .io_enq_last(NothingFilter_1_io_enq_last),
    .io_deq_ready(NothingFilter_1_io_deq_ready),
    .io_deq_valid(NothingFilter_1_io_deq_valid),
    .io_deq_bits(NothingFilter_1_io_deq_bits),
    .io_deq_user(NothingFilter_1_io_deq_user),
    .io_deq_last(NothingFilter_1_io_deq_last)
  );
  NothingFilter NothingFilter_2 ( // @[ChiselImProc.scala 469:16]
    .clock(NothingFilter_2_clock),
    .reset(NothingFilter_2_reset),
    .io_enq_ready(NothingFilter_2_io_enq_ready),
    .io_enq_valid(NothingFilter_2_io_enq_valid),
    .io_enq_bits(NothingFilter_2_io_enq_bits),
    .io_enq_user(NothingFilter_2_io_enq_user),
    .io_enq_last(NothingFilter_2_io_enq_last),
    .io_deq_ready(NothingFilter_2_io_deq_ready),
    .io_deq_valid(NothingFilter_2_io_deq_valid),
    .io_deq_bits(NothingFilter_2_io_deq_bits),
    .io_deq_user(NothingFilter_2_io_deq_user),
    .io_deq_last(NothingFilter_2_io_deq_last)
  );
  NothingFilter NothingFilter_3 ( // @[ChiselImProc.scala 472:16]
    .clock(NothingFilter_3_clock),
    .reset(NothingFilter_3_reset),
    .io_enq_ready(NothingFilter_3_io_enq_ready),
    .io_enq_valid(NothingFilter_3_io_enq_valid),
    .io_enq_bits(NothingFilter_3_io_enq_bits),
    .io_enq_user(NothingFilter_3_io_enq_user),
    .io_enq_last(NothingFilter_3_io_enq_last),
    .io_deq_ready(NothingFilter_3_io_deq_ready),
    .io_deq_valid(NothingFilter_3_io_deq_valid),
    .io_deq_bits(NothingFilter_3_io_deq_bits),
    .io_deq_user(NothingFilter_3_io_deq_user),
    .io_deq_last(NothingFilter_3_io_deq_last)
  );
  Gray2RGBFilter Gray2RGBFilter ( // @[ChiselImProc.scala 474:16]
    .clock(Gray2RGBFilter_clock),
    .reset(Gray2RGBFilter_reset),
    .io_enq_ready(Gray2RGBFilter_io_enq_ready),
    .io_enq_valid(Gray2RGBFilter_io_enq_valid),
    .io_enq_bits(Gray2RGBFilter_io_enq_bits),
    .io_enq_user(Gray2RGBFilter_io_enq_user),
    .io_enq_last(Gray2RGBFilter_io_enq_last),
    .io_deq_ready(Gray2RGBFilter_io_deq_ready),
    .io_deq_valid(Gray2RGBFilter_io_deq_valid),
    .io_deq_bits(Gray2RGBFilter_io_deq_bits),
    .io_deq_user(Gray2RGBFilter_io_deq_user),
    .io_deq_last(Gray2RGBFilter_io_deq_last)
  );
  assign io_enq_ready = RGB2GrayFilter_io_enq_ready; // @[ChiselImProc.scala 485:12]
  assign io_deq_valid = Gray2RGBFilter_io_deq_valid; // @[ChiselImProc.scala 487:12]
  assign io_deq_bits = Gray2RGBFilter_io_deq_bits; // @[ChiselImProc.scala 487:12]
  assign io_deq_user = Gray2RGBFilter_io_deq_user; // @[ChiselImProc.scala 487:12]
  assign io_deq_last = Gray2RGBFilter_io_deq_last; // @[ChiselImProc.scala 487:12]
  assign io_dport = 32'h0; // @[ChiselImProc.scala 505:14]
  assign io_dport2 = 32'h0; // @[ChiselImProc.scala 506:15]
  assign RGB2GrayFilter_clock = clock;
  assign RGB2GrayFilter_reset = reset;
  assign RGB2GrayFilter_io_enq_valid = io_enq_valid; // @[ChiselImProc.scala 485:12]
  assign RGB2GrayFilter_io_enq_bits = io_enq_bits; // @[ChiselImProc.scala 485:12]
  assign RGB2GrayFilter_io_enq_user = io_enq_user; // @[ChiselImProc.scala 485:12]
  assign RGB2GrayFilter_io_enq_last = io_enq_last; // @[ChiselImProc.scala 485:12]
  assign RGB2GrayFilter_io_deq_ready = GaussianBlurFilter_io_enq_ready; // @[ChiselImProc.scala 482:30]
  assign GaussianBlurFilter_clock = clock;
  assign GaussianBlurFilter_reset = reset;
  assign GaussianBlurFilter_io_enq_valid = RGB2GrayFilter_io_deq_valid; // @[ChiselImProc.scala 482:30]
  assign GaussianBlurFilter_io_enq_bits = RGB2GrayFilter_io_deq_bits[7:0]; // @[ChiselImProc.scala 482:30]
  assign GaussianBlurFilter_io_enq_user = RGB2GrayFilter_io_deq_user; // @[ChiselImProc.scala 482:30]
  assign GaussianBlurFilter_io_enq_last = RGB2GrayFilter_io_deq_last; // @[ChiselImProc.scala 482:30]
  assign GaussianBlurFilter_io_deq_ready = NothingFilter_io_enq_ready; // @[ChiselImProc.scala 482:30]
  assign NothingFilter_clock = clock;
  assign NothingFilter_reset = reset;
  assign NothingFilter_io_enq_valid = GaussianBlurFilter_io_deq_valid; // @[ChiselImProc.scala 482:30]
  assign NothingFilter_io_enq_bits = GaussianBlurFilter_io_deq_bits; // @[ChiselImProc.scala 482:30]
  assign NothingFilter_io_enq_user = GaussianBlurFilter_io_deq_user; // @[ChiselImProc.scala 482:30]
  assign NothingFilter_io_enq_last = GaussianBlurFilter_io_deq_last; // @[ChiselImProc.scala 482:30]
  assign NothingFilter_io_deq_ready = NothingFilter_1_io_enq_ready; // @[ChiselImProc.scala 482:30]
  assign NothingFilter_1_clock = clock;
  assign NothingFilter_1_reset = reset;
  assign NothingFilter_1_io_enq_valid = NothingFilter_io_deq_valid; // @[ChiselImProc.scala 482:30]
  assign NothingFilter_1_io_enq_bits = NothingFilter_io_deq_bits; // @[ChiselImProc.scala 482:30]
  assign NothingFilter_1_io_enq_user = NothingFilter_io_deq_user; // @[ChiselImProc.scala 482:30]
  assign NothingFilter_1_io_enq_last = NothingFilter_io_deq_last; // @[ChiselImProc.scala 482:30]
  assign NothingFilter_1_io_deq_ready = NothingFilter_2_io_enq_ready; // @[ChiselImProc.scala 482:30]
  assign NothingFilter_2_clock = clock;
  assign NothingFilter_2_reset = reset;
  assign NothingFilter_2_io_enq_valid = NothingFilter_1_io_deq_valid; // @[ChiselImProc.scala 482:30]
  assign NothingFilter_2_io_enq_bits = NothingFilter_1_io_deq_bits; // @[ChiselImProc.scala 482:30]
  assign NothingFilter_2_io_enq_user = NothingFilter_1_io_deq_user; // @[ChiselImProc.scala 482:30]
  assign NothingFilter_2_io_enq_last = NothingFilter_1_io_deq_last; // @[ChiselImProc.scala 482:30]
  assign NothingFilter_2_io_deq_ready = NothingFilter_3_io_enq_ready; // @[ChiselImProc.scala 482:30]
  assign NothingFilter_3_clock = clock;
  assign NothingFilter_3_reset = reset;
  assign NothingFilter_3_io_enq_valid = NothingFilter_2_io_deq_valid; // @[ChiselImProc.scala 482:30]
  assign NothingFilter_3_io_enq_bits = NothingFilter_2_io_deq_bits; // @[ChiselImProc.scala 482:30]
  assign NothingFilter_3_io_enq_user = NothingFilter_2_io_deq_user; // @[ChiselImProc.scala 482:30]
  assign NothingFilter_3_io_enq_last = NothingFilter_2_io_deq_last; // @[ChiselImProc.scala 482:30]
  assign NothingFilter_3_io_deq_ready = Gray2RGBFilter_io_enq_ready; // @[ChiselImProc.scala 482:30]
  assign Gray2RGBFilter_clock = clock;
  assign Gray2RGBFilter_reset = reset;
  assign Gray2RGBFilter_io_enq_valid = NothingFilter_3_io_deq_valid; // @[ChiselImProc.scala 482:30]
  assign Gray2RGBFilter_io_enq_bits = {{16'd0}, NothingFilter_3_io_deq_bits}; // @[ChiselImProc.scala 482:30]
  assign Gray2RGBFilter_io_enq_user = NothingFilter_3_io_deq_user; // @[ChiselImProc.scala 482:30]
  assign Gray2RGBFilter_io_enq_last = NothingFilter_3_io_deq_last; // @[ChiselImProc.scala 482:30]
  assign Gray2RGBFilter_io_deq_ready = io_deq_ready; // @[ChiselImProc.scala 487:12]
endmodule

module SqrtExtractionUInt(
  input         clock,
  input         reset,
  input  [15:0] io_z,
  output [7:0]  io_q
);
  wire [16:0] zj_7 = {1'h0,io_z[15:14],14'h0}; // @[Cat.scala 29:58]
  wire [2:0] _T_5 = zj_7[16:14] - 3'h1; // @[Sqrt.scala 54:77]
  wire [16:0] rj_7 = {_T_5,14'h0}; // @[Cat.scala 29:58]
  wire  qSub_7 = ~rj_7[16]; // @[Sqrt.scala 55:27]
  wire [4:0] _T_11 = {rj_7[16:14],io_z[13:12]}; // @[Cat.scala 29:58]
  wire [16:0] _GEN_7 = {_T_11, 12'h0}; // @[Sqrt.scala 59:77]
  wire [19:0] _T_12 = {{3'd0}, _GEN_7}; // @[Sqrt.scala 59:77]
  wire [4:0] _T_15 = {zj_7[16:14],io_z[13:12]}; // @[Cat.scala 29:58]
  wire [16:0] _GEN_8 = {_T_15, 12'h0}; // @[Sqrt.scala 61:77]
  wire [19:0] _T_16 = {{3'd0}, _GEN_8}; // @[Sqrt.scala 61:77]
  wire [19:0] _GEN_0 = qSub_7 ? _T_12 : _T_16; // @[Sqrt.scala 58:26]
  wire [16:0] zj_6 = _GEN_0[16:0]; // @[Sqrt.scala 47:19 Sqrt.scala 59:19 Sqrt.scala 61:19]
  wire [2:0] _T_20 = {qSub_7,2'h1}; // @[Cat.scala 29:58]
  wire [4:0] _GEN_9 = {{2'd0}, _T_20}; // @[Sqrt.scala 64:45]
  wire [4:0] _T_22 = zj_6[16:12] - _GEN_9; // @[Sqrt.scala 64:45]
  wire [16:0] _GEN_10 = {_T_22, 12'h0}; // @[Sqrt.scala 64:77]
  wire [19:0] _T_23 = {{3'd0}, _GEN_10}; // @[Sqrt.scala 64:77]
  wire [16:0] rj_6 = _T_23[16:0]; // @[Sqrt.scala 48:19 Sqrt.scala 64:15]
  wire  qSub_6 = ~rj_6[16]; // @[Sqrt.scala 65:20]
  wire [5:0] _T_28 = {rj_6[15:12],io_z[11:10]}; // @[Cat.scala 29:58]
  wire [15:0] _GEN_11 = {_T_28, 10'h0}; // @[Sqrt.scala 59:77]
  wire [20:0] _T_29 = {{5'd0}, _GEN_11}; // @[Sqrt.scala 59:77]
  wire [5:0] _T_32 = {zj_6[15:12],io_z[11:10]}; // @[Cat.scala 29:58]
  wire [15:0] _GEN_12 = {_T_32, 10'h0}; // @[Sqrt.scala 61:77]
  wire [20:0] _T_33 = {{5'd0}, _GEN_12}; // @[Sqrt.scala 61:77]
  wire [20:0] _GEN_1 = qSub_6 ? _T_29 : _T_33; // @[Sqrt.scala 58:26]
  wire [16:0] zj_5 = _GEN_1[16:0]; // @[Sqrt.scala 47:19 Sqrt.scala 59:19 Sqrt.scala 61:19]
  wire [3:0] _T_38 = {qSub_7,qSub_6,2'h1}; // @[Cat.scala 29:58]
  wire [5:0] _GEN_13 = {{2'd0}, _T_38}; // @[Sqrt.scala 64:45]
  wire [5:0] _T_40 = zj_5[15:10] - _GEN_13; // @[Sqrt.scala 64:45]
  wire [15:0] _GEN_14 = {_T_40, 10'h0}; // @[Sqrt.scala 64:77]
  wire [20:0] _T_41 = {{5'd0}, _GEN_14}; // @[Sqrt.scala 64:77]
  wire [16:0] rj_5 = _T_41[16:0]; // @[Sqrt.scala 48:19 Sqrt.scala 64:15]
  wire  qSub_5 = ~rj_5[15]; // @[Sqrt.scala 65:20]
  wire [6:0] _T_46 = {rj_5[14:10],io_z[9:8]}; // @[Cat.scala 29:58]
  wire [14:0] _GEN_15 = {_T_46, 8'h0}; // @[Sqrt.scala 59:77]
  wire [21:0] _T_47 = {{7'd0}, _GEN_15}; // @[Sqrt.scala 59:77]
  wire [6:0] _T_50 = {zj_5[14:10],io_z[9:8]}; // @[Cat.scala 29:58]
  wire [14:0] _GEN_16 = {_T_50, 8'h0}; // @[Sqrt.scala 61:77]
  wire [21:0] _T_51 = {{7'd0}, _GEN_16}; // @[Sqrt.scala 61:77]
  wire [21:0] _GEN_2 = qSub_5 ? _T_47 : _T_51; // @[Sqrt.scala 58:26]
  wire [16:0] zj_4 = _GEN_2[16:0]; // @[Sqrt.scala 47:19 Sqrt.scala 59:19 Sqrt.scala 61:19]
  wire [4:0] _T_57 = {qSub_7,qSub_6,qSub_5,2'h1}; // @[Cat.scala 29:58]
  wire [6:0] _GEN_17 = {{2'd0}, _T_57}; // @[Sqrt.scala 64:45]
  wire [6:0] _T_59 = zj_4[14:8] - _GEN_17; // @[Sqrt.scala 64:45]
  wire [14:0] _GEN_18 = {_T_59, 8'h0}; // @[Sqrt.scala 64:77]
  wire [21:0] _T_60 = {{7'd0}, _GEN_18}; // @[Sqrt.scala 64:77]
  wire [16:0] rj_4 = _T_60[16:0]; // @[Sqrt.scala 48:19 Sqrt.scala 64:15]
  wire  qSub_4 = ~rj_4[14]; // @[Sqrt.scala 65:20]
  wire [7:0] _T_65 = {rj_4[13:8],io_z[7:6]}; // @[Cat.scala 29:58]
  wire [13:0] _GEN_19 = {_T_65, 6'h0}; // @[Sqrt.scala 59:77]
  wire [14:0] _T_66 = {{1'd0}, _GEN_19}; // @[Sqrt.scala 59:77]
  wire [7:0] _T_69 = {zj_4[13:8],io_z[7:6]}; // @[Cat.scala 29:58]
  wire [13:0] _GEN_20 = {_T_69, 6'h0}; // @[Sqrt.scala 61:77]
  wire [14:0] _T_70 = {{1'd0}, _GEN_20}; // @[Sqrt.scala 61:77]
  wire [14:0] _GEN_3 = qSub_4 ? _T_66 : _T_70; // @[Sqrt.scala 58:26]
  wire [16:0] zj_3 = {{2'd0}, _GEN_3}; // @[Sqrt.scala 47:19 Sqrt.scala 59:19 Sqrt.scala 61:19]
  wire [3:0] _T_76 = {qSub_7,qSub_6,qSub_5,qSub_4}; // @[Sqrt.scala 64:58]
  wire [5:0] _T_77 = {qSub_7,qSub_6,qSub_5,qSub_4,2'h1}; // @[Cat.scala 29:58]
  wire [7:0] _GEN_21 = {{2'd0}, _T_77}; // @[Sqrt.scala 64:45]
  wire [7:0] _T_79 = zj_3[13:6] - _GEN_21; // @[Sqrt.scala 64:45]
  wire [13:0] _GEN_22 = {_T_79, 6'h0}; // @[Sqrt.scala 64:77]
  wire [14:0] _T_80 = {{1'd0}, _GEN_22}; // @[Sqrt.scala 64:77]
  wire [16:0] rj_3 = {{2'd0}, _T_80}; // @[Sqrt.scala 48:19 Sqrt.scala 64:15]
  wire  qSub_3 = ~rj_3[13]; // @[Sqrt.scala 65:20]
  wire [8:0] _T_85 = {rj_3[12:6],io_z[5:4]}; // @[Cat.scala 29:58]
  wire [12:0] _GEN_23 = {_T_85, 4'h0}; // @[Sqrt.scala 59:77]
  wire [15:0] _T_86 = {{3'd0}, _GEN_23}; // @[Sqrt.scala 59:77]
  wire [8:0] _T_89 = {zj_3[12:6],io_z[5:4]}; // @[Cat.scala 29:58]
  wire [12:0] _GEN_24 = {_T_89, 4'h0}; // @[Sqrt.scala 61:77]
  wire [15:0] _T_90 = {{3'd0}, _GEN_24}; // @[Sqrt.scala 61:77]
  wire [15:0] _GEN_4 = qSub_3 ? _T_86 : _T_90; // @[Sqrt.scala 58:26]
  wire [16:0] zj_2 = {{1'd0}, _GEN_4}; // @[Sqrt.scala 47:19 Sqrt.scala 59:19 Sqrt.scala 61:19]
  wire [6:0] _T_98 = {qSub_7,qSub_6,qSub_5,qSub_4,qSub_3,2'h1}; // @[Cat.scala 29:58]
  wire [8:0] _GEN_25 = {{2'd0}, _T_98}; // @[Sqrt.scala 64:45]
  wire [8:0] _T_100 = zj_2[12:4] - _GEN_25; // @[Sqrt.scala 64:45]
  wire [12:0] _GEN_26 = {_T_100, 4'h0}; // @[Sqrt.scala 64:77]
  wire [15:0] _T_101 = {{3'd0}, _GEN_26}; // @[Sqrt.scala 64:77]
  wire [16:0] rj_2 = {{1'd0}, _T_101}; // @[Sqrt.scala 48:19 Sqrt.scala 64:15]
  wire  qSub_2 = ~rj_2[12]; // @[Sqrt.scala 65:20]
  wire [9:0] _T_106 = {rj_2[11:4],io_z[3:2]}; // @[Cat.scala 29:58]
  wire [11:0] _GEN_27 = {_T_106, 2'h0}; // @[Sqrt.scala 59:77]
  wire [12:0] _T_107 = {{1'd0}, _GEN_27}; // @[Sqrt.scala 59:77]
  wire [9:0] _T_110 = {zj_2[11:4],io_z[3:2]}; // @[Cat.scala 29:58]
  wire [11:0] _GEN_28 = {_T_110, 2'h0}; // @[Sqrt.scala 61:77]
  wire [12:0] _T_111 = {{1'd0}, _GEN_28}; // @[Sqrt.scala 61:77]
  wire [12:0] _GEN_5 = qSub_2 ? _T_107 : _T_111; // @[Sqrt.scala 58:26]
  wire [16:0] zj_1 = {{4'd0}, _GEN_5}; // @[Sqrt.scala 47:19 Sqrt.scala 59:19 Sqrt.scala 61:19]
  wire [7:0] _T_120 = {qSub_7,qSub_6,qSub_5,qSub_4,qSub_3,qSub_2,2'h1}; // @[Cat.scala 29:58]
  wire [9:0] _GEN_29 = {{2'd0}, _T_120}; // @[Sqrt.scala 64:45]
  wire [9:0] _T_122 = zj_1[11:2] - _GEN_29; // @[Sqrt.scala 64:45]
  wire [11:0] _GEN_30 = {_T_122, 2'h0}; // @[Sqrt.scala 64:77]
  wire [12:0] _T_123 = {{1'd0}, _GEN_30}; // @[Sqrt.scala 64:77]
  wire [16:0] rj_1 = {{4'd0}, _T_123}; // @[Sqrt.scala 48:19 Sqrt.scala 64:15]
  wire  qSub_1 = ~rj_1[11]; // @[Sqrt.scala 65:20]
  wire [10:0] _T_128 = {rj_1[10:2],io_z[1:0]}; // @[Cat.scala 29:58]
  wire [11:0] _T_129 = {{1'd0}, _T_128}; // @[Sqrt.scala 59:77]
  wire [10:0] _T_132 = {zj_1[10:2],io_z[1:0]}; // @[Cat.scala 29:58]
  wire [11:0] _T_133 = {{1'd0}, _T_132}; // @[Sqrt.scala 61:77]
  wire [11:0] _GEN_6 = qSub_1 ? _T_129 : _T_133; // @[Sqrt.scala 58:26]
  wire [16:0] zj_0 = {{5'd0}, _GEN_6}; // @[Sqrt.scala 47:19 Sqrt.scala 59:19 Sqrt.scala 61:19]
  wire [8:0] _T_143 = {qSub_7,qSub_6,qSub_5,qSub_4,qSub_3,qSub_2,qSub_1,2'h1}; // @[Cat.scala 29:58]
  wire [10:0] _GEN_31 = {{2'd0}, _T_143}; // @[Sqrt.scala 64:45]
  wire [10:0] _T_145 = zj_0[10:0] - _GEN_31; // @[Sqrt.scala 64:45]
  wire [11:0] _T_146 = {{1'd0}, _T_145}; // @[Sqrt.scala 64:77]
  wire [16:0] rj_0 = {{5'd0}, _T_146}; // @[Sqrt.scala 48:19 Sqrt.scala 64:15]
  wire  qSub_0 = ~rj_0[10]; // @[Sqrt.scala 65:20]
  wire [3:0] _T_151 = {qSub_3,qSub_2,qSub_1,qSub_0}; // @[Sqrt.scala 68:18]
  assign io_q = {_T_76,_T_151}; // @[Sqrt.scala 68:10]
endmodule
